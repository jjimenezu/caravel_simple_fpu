magic
tech sky130A
magscale 1 2
timestamp 1733387643
<< obsli1 >>
rect 1104 2159 135148 136017
<< obsm1 >>
rect 198 1232 136054 136264
<< metal2 >>
rect 3514 137670 3570 138470
rect 8482 137670 8538 138470
rect 13450 137670 13506 138470
rect 18418 137670 18474 138470
rect 23386 137670 23442 138470
rect 28354 137670 28410 138470
rect 33322 137670 33378 138470
rect 38290 137670 38346 138470
rect 43258 137670 43314 138470
rect 48226 137670 48282 138470
rect 53194 137670 53250 138470
rect 58162 137670 58218 138470
rect 63130 137670 63186 138470
rect 68098 137670 68154 138470
rect 73066 137670 73122 138470
rect 78034 137670 78090 138470
rect 83002 137670 83058 138470
rect 87970 137670 88026 138470
rect 92938 137670 92994 138470
rect 97906 137670 97962 138470
rect 102874 137670 102930 138470
rect 107842 137670 107898 138470
rect 112810 137670 112866 138470
rect 117778 137670 117834 138470
rect 122746 137670 122802 138470
rect 127714 137670 127770 138470
rect 132682 137670 132738 138470
rect 202 0 258 800
rect 478 0 534 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1582 0 1638 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2410 0 2466 800
rect 2686 0 2742 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 4066 0 4122 800
rect 4342 0 4398 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5722 0 5778 800
rect 5998 0 6054 800
rect 6274 0 6330 800
rect 6550 0 6606 800
rect 6826 0 6882 800
rect 7102 0 7158 800
rect 7378 0 7434 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8482 0 8538 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10138 0 10194 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 10966 0 11022 800
rect 11242 0 11298 800
rect 11518 0 11574 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27250 0 27306 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29458 0 29514 800
rect 29734 0 29790 800
rect 30010 0 30066 800
rect 30286 0 30342 800
rect 30562 0 30618 800
rect 30838 0 30894 800
rect 31114 0 31170 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32770 0 32826 800
rect 33046 0 33102 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33874 0 33930 800
rect 34150 0 34206 800
rect 34426 0 34482 800
rect 34702 0 34758 800
rect 34978 0 35034 800
rect 35254 0 35310 800
rect 35530 0 35586 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36634 0 36690 800
rect 36910 0 36966 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39394 0 39450 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40774 0 40830 800
rect 41050 0 41106 800
rect 41326 0 41382 800
rect 41602 0 41658 800
rect 41878 0 41934 800
rect 42154 0 42210 800
rect 42430 0 42486 800
rect 42706 0 42762 800
rect 42982 0 43038 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44362 0 44418 800
rect 44638 0 44694 800
rect 44914 0 44970 800
rect 45190 0 45246 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 46018 0 46074 800
rect 46294 0 46350 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47122 0 47178 800
rect 47398 0 47454 800
rect 47674 0 47730 800
rect 47950 0 48006 800
rect 48226 0 48282 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49882 0 49938 800
rect 50158 0 50214 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51262 0 51318 800
rect 51538 0 51594 800
rect 51814 0 51870 800
rect 52090 0 52146 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53194 0 53250 800
rect 53470 0 53526 800
rect 53746 0 53802 800
rect 54022 0 54078 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54850 0 54906 800
rect 55126 0 55182 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 55954 0 56010 800
rect 56230 0 56286 800
rect 56506 0 56562 800
rect 56782 0 56838 800
rect 57058 0 57114 800
rect 57334 0 57390 800
rect 57610 0 57666 800
rect 57886 0 57942 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58714 0 58770 800
rect 58990 0 59046 800
rect 59266 0 59322 800
rect 59542 0 59598 800
rect 59818 0 59874 800
rect 60094 0 60150 800
rect 60370 0 60426 800
rect 60646 0 60702 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61474 0 61530 800
rect 61750 0 61806 800
rect 62026 0 62082 800
rect 62302 0 62358 800
rect 62578 0 62634 800
rect 62854 0 62910 800
rect 63130 0 63186 800
rect 63406 0 63462 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64234 0 64290 800
rect 64510 0 64566 800
rect 64786 0 64842 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66442 0 66498 800
rect 66718 0 66774 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67546 0 67602 800
rect 67822 0 67878 800
rect 68098 0 68154 800
rect 68374 0 68430 800
rect 68650 0 68706 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70306 0 70362 800
rect 70582 0 70638 800
rect 70858 0 70914 800
rect 71134 0 71190 800
rect 71410 0 71466 800
rect 71686 0 71742 800
rect 71962 0 72018 800
rect 72238 0 72294 800
rect 72514 0 72570 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73342 0 73398 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74170 0 74226 800
rect 74446 0 74502 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75550 0 75606 800
rect 75826 0 75882 800
rect 76102 0 76158 800
rect 76378 0 76434 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77206 0 77262 800
rect 77482 0 77538 800
rect 77758 0 77814 800
rect 78034 0 78090 800
rect 78310 0 78366 800
rect 78586 0 78642 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79690 0 79746 800
rect 79966 0 80022 800
rect 80242 0 80298 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 81070 0 81126 800
rect 81346 0 81402 800
rect 81622 0 81678 800
rect 81898 0 81954 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82726 0 82782 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83554 0 83610 800
rect 83830 0 83886 800
rect 84106 0 84162 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84934 0 84990 800
rect 85210 0 85266 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86314 0 86370 800
rect 86590 0 86646 800
rect 86866 0 86922 800
rect 87142 0 87198 800
rect 87418 0 87474 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 89074 0 89130 800
rect 89350 0 89406 800
rect 89626 0 89682 800
rect 89902 0 89958 800
rect 90178 0 90234 800
rect 90454 0 90510 800
rect 90730 0 90786 800
rect 91006 0 91062 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91834 0 91890 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92662 0 92718 800
rect 92938 0 92994 800
rect 93214 0 93270 800
rect 93490 0 93546 800
rect 93766 0 93822 800
rect 94042 0 94098 800
rect 94318 0 94374 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95698 0 95754 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97354 0 97410 800
rect 97630 0 97686 800
rect 97906 0 97962 800
rect 98182 0 98238 800
rect 98458 0 98514 800
rect 98734 0 98790 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99562 0 99618 800
rect 99838 0 99894 800
rect 100114 0 100170 800
rect 100390 0 100446 800
rect 100666 0 100722 800
rect 100942 0 100998 800
rect 101218 0 101274 800
rect 101494 0 101550 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102322 0 102378 800
rect 102598 0 102654 800
rect 102874 0 102930 800
rect 103150 0 103206 800
rect 103426 0 103482 800
rect 103702 0 103758 800
rect 103978 0 104034 800
rect 104254 0 104310 800
rect 104530 0 104586 800
rect 104806 0 104862 800
rect 105082 0 105138 800
rect 105358 0 105414 800
rect 105634 0 105690 800
rect 105910 0 105966 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106738 0 106794 800
rect 107014 0 107070 800
rect 107290 0 107346 800
rect 107566 0 107622 800
rect 107842 0 107898 800
rect 108118 0 108174 800
rect 108394 0 108450 800
rect 108670 0 108726 800
rect 108946 0 109002 800
rect 109222 0 109278 800
rect 109498 0 109554 800
rect 109774 0 109830 800
rect 110050 0 110106 800
rect 110326 0 110382 800
rect 110602 0 110658 800
rect 110878 0 110934 800
rect 111154 0 111210 800
rect 111430 0 111486 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112258 0 112314 800
rect 112534 0 112590 800
rect 112810 0 112866 800
rect 113086 0 113142 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 113914 0 113970 800
rect 114190 0 114246 800
rect 114466 0 114522 800
rect 114742 0 114798 800
rect 115018 0 115074 800
rect 115294 0 115350 800
rect 115570 0 115626 800
rect 115846 0 115902 800
rect 116122 0 116178 800
rect 116398 0 116454 800
rect 116674 0 116730 800
rect 116950 0 117006 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117778 0 117834 800
rect 118054 0 118110 800
rect 118330 0 118386 800
rect 118606 0 118662 800
rect 118882 0 118938 800
rect 119158 0 119214 800
rect 119434 0 119490 800
rect 119710 0 119766 800
rect 119986 0 120042 800
rect 120262 0 120318 800
rect 120538 0 120594 800
rect 120814 0 120870 800
rect 121090 0 121146 800
rect 121366 0 121422 800
rect 121642 0 121698 800
rect 121918 0 121974 800
rect 122194 0 122250 800
rect 122470 0 122526 800
rect 122746 0 122802 800
rect 123022 0 123078 800
rect 123298 0 123354 800
rect 123574 0 123630 800
rect 123850 0 123906 800
rect 124126 0 124182 800
rect 124402 0 124458 800
rect 124678 0 124734 800
rect 124954 0 125010 800
rect 125230 0 125286 800
rect 125506 0 125562 800
rect 125782 0 125838 800
rect 126058 0 126114 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126886 0 126942 800
rect 127162 0 127218 800
rect 127438 0 127494 800
rect 127714 0 127770 800
rect 127990 0 128046 800
rect 128266 0 128322 800
rect 128542 0 128598 800
rect 128818 0 128874 800
rect 129094 0 129150 800
rect 129370 0 129426 800
rect 129646 0 129702 800
rect 129922 0 129978 800
rect 130198 0 130254 800
rect 130474 0 130530 800
rect 130750 0 130806 800
rect 131026 0 131082 800
rect 131302 0 131358 800
rect 131578 0 131634 800
rect 131854 0 131910 800
rect 132130 0 132186 800
rect 132406 0 132462 800
rect 132682 0 132738 800
rect 132958 0 133014 800
rect 133234 0 133290 800
rect 133510 0 133566 800
rect 133786 0 133842 800
rect 134062 0 134118 800
rect 134338 0 134394 800
rect 134614 0 134670 800
rect 134890 0 134946 800
rect 135166 0 135222 800
rect 135442 0 135498 800
rect 135718 0 135774 800
rect 135994 0 136050 800
<< obsm2 >>
rect 204 137614 3458 137670
rect 3626 137614 8426 137670
rect 8594 137614 13394 137670
rect 13562 137614 18362 137670
rect 18530 137614 23330 137670
rect 23498 137614 28298 137670
rect 28466 137614 33266 137670
rect 33434 137614 38234 137670
rect 38402 137614 43202 137670
rect 43370 137614 48170 137670
rect 48338 137614 53138 137670
rect 53306 137614 58106 137670
rect 58274 137614 63074 137670
rect 63242 137614 68042 137670
rect 68210 137614 73010 137670
rect 73178 137614 77978 137670
rect 78146 137614 82946 137670
rect 83114 137614 87914 137670
rect 88082 137614 92882 137670
rect 93050 137614 97850 137670
rect 98018 137614 102818 137670
rect 102986 137614 107786 137670
rect 107954 137614 112754 137670
rect 112922 137614 117722 137670
rect 117890 137614 122690 137670
rect 122858 137614 127658 137670
rect 127826 137614 132626 137670
rect 132794 137614 136048 137670
rect 204 856 136048 137614
rect 314 800 422 856
rect 590 800 698 856
rect 866 800 974 856
rect 1142 800 1250 856
rect 1418 800 1526 856
rect 1694 800 1802 856
rect 1970 800 2078 856
rect 2246 800 2354 856
rect 2522 800 2630 856
rect 2798 800 2906 856
rect 3074 800 3182 856
rect 3350 800 3458 856
rect 3626 800 3734 856
rect 3902 800 4010 856
rect 4178 800 4286 856
rect 4454 800 4562 856
rect 4730 800 4838 856
rect 5006 800 5114 856
rect 5282 800 5390 856
rect 5558 800 5666 856
rect 5834 800 5942 856
rect 6110 800 6218 856
rect 6386 800 6494 856
rect 6662 800 6770 856
rect 6938 800 7046 856
rect 7214 800 7322 856
rect 7490 800 7598 856
rect 7766 800 7874 856
rect 8042 800 8150 856
rect 8318 800 8426 856
rect 8594 800 8702 856
rect 8870 800 8978 856
rect 9146 800 9254 856
rect 9422 800 9530 856
rect 9698 800 9806 856
rect 9974 800 10082 856
rect 10250 800 10358 856
rect 10526 800 10634 856
rect 10802 800 10910 856
rect 11078 800 11186 856
rect 11354 800 11462 856
rect 11630 800 11738 856
rect 11906 800 12014 856
rect 12182 800 12290 856
rect 12458 800 12566 856
rect 12734 800 12842 856
rect 13010 800 13118 856
rect 13286 800 13394 856
rect 13562 800 13670 856
rect 13838 800 13946 856
rect 14114 800 14222 856
rect 14390 800 14498 856
rect 14666 800 14774 856
rect 14942 800 15050 856
rect 15218 800 15326 856
rect 15494 800 15602 856
rect 15770 800 15878 856
rect 16046 800 16154 856
rect 16322 800 16430 856
rect 16598 800 16706 856
rect 16874 800 16982 856
rect 17150 800 17258 856
rect 17426 800 17534 856
rect 17702 800 17810 856
rect 17978 800 18086 856
rect 18254 800 18362 856
rect 18530 800 18638 856
rect 18806 800 18914 856
rect 19082 800 19190 856
rect 19358 800 19466 856
rect 19634 800 19742 856
rect 19910 800 20018 856
rect 20186 800 20294 856
rect 20462 800 20570 856
rect 20738 800 20846 856
rect 21014 800 21122 856
rect 21290 800 21398 856
rect 21566 800 21674 856
rect 21842 800 21950 856
rect 22118 800 22226 856
rect 22394 800 22502 856
rect 22670 800 22778 856
rect 22946 800 23054 856
rect 23222 800 23330 856
rect 23498 800 23606 856
rect 23774 800 23882 856
rect 24050 800 24158 856
rect 24326 800 24434 856
rect 24602 800 24710 856
rect 24878 800 24986 856
rect 25154 800 25262 856
rect 25430 800 25538 856
rect 25706 800 25814 856
rect 25982 800 26090 856
rect 26258 800 26366 856
rect 26534 800 26642 856
rect 26810 800 26918 856
rect 27086 800 27194 856
rect 27362 800 27470 856
rect 27638 800 27746 856
rect 27914 800 28022 856
rect 28190 800 28298 856
rect 28466 800 28574 856
rect 28742 800 28850 856
rect 29018 800 29126 856
rect 29294 800 29402 856
rect 29570 800 29678 856
rect 29846 800 29954 856
rect 30122 800 30230 856
rect 30398 800 30506 856
rect 30674 800 30782 856
rect 30950 800 31058 856
rect 31226 800 31334 856
rect 31502 800 31610 856
rect 31778 800 31886 856
rect 32054 800 32162 856
rect 32330 800 32438 856
rect 32606 800 32714 856
rect 32882 800 32990 856
rect 33158 800 33266 856
rect 33434 800 33542 856
rect 33710 800 33818 856
rect 33986 800 34094 856
rect 34262 800 34370 856
rect 34538 800 34646 856
rect 34814 800 34922 856
rect 35090 800 35198 856
rect 35366 800 35474 856
rect 35642 800 35750 856
rect 35918 800 36026 856
rect 36194 800 36302 856
rect 36470 800 36578 856
rect 36746 800 36854 856
rect 37022 800 37130 856
rect 37298 800 37406 856
rect 37574 800 37682 856
rect 37850 800 37958 856
rect 38126 800 38234 856
rect 38402 800 38510 856
rect 38678 800 38786 856
rect 38954 800 39062 856
rect 39230 800 39338 856
rect 39506 800 39614 856
rect 39782 800 39890 856
rect 40058 800 40166 856
rect 40334 800 40442 856
rect 40610 800 40718 856
rect 40886 800 40994 856
rect 41162 800 41270 856
rect 41438 800 41546 856
rect 41714 800 41822 856
rect 41990 800 42098 856
rect 42266 800 42374 856
rect 42542 800 42650 856
rect 42818 800 42926 856
rect 43094 800 43202 856
rect 43370 800 43478 856
rect 43646 800 43754 856
rect 43922 800 44030 856
rect 44198 800 44306 856
rect 44474 800 44582 856
rect 44750 800 44858 856
rect 45026 800 45134 856
rect 45302 800 45410 856
rect 45578 800 45686 856
rect 45854 800 45962 856
rect 46130 800 46238 856
rect 46406 800 46514 856
rect 46682 800 46790 856
rect 46958 800 47066 856
rect 47234 800 47342 856
rect 47510 800 47618 856
rect 47786 800 47894 856
rect 48062 800 48170 856
rect 48338 800 48446 856
rect 48614 800 48722 856
rect 48890 800 48998 856
rect 49166 800 49274 856
rect 49442 800 49550 856
rect 49718 800 49826 856
rect 49994 800 50102 856
rect 50270 800 50378 856
rect 50546 800 50654 856
rect 50822 800 50930 856
rect 51098 800 51206 856
rect 51374 800 51482 856
rect 51650 800 51758 856
rect 51926 800 52034 856
rect 52202 800 52310 856
rect 52478 800 52586 856
rect 52754 800 52862 856
rect 53030 800 53138 856
rect 53306 800 53414 856
rect 53582 800 53690 856
rect 53858 800 53966 856
rect 54134 800 54242 856
rect 54410 800 54518 856
rect 54686 800 54794 856
rect 54962 800 55070 856
rect 55238 800 55346 856
rect 55514 800 55622 856
rect 55790 800 55898 856
rect 56066 800 56174 856
rect 56342 800 56450 856
rect 56618 800 56726 856
rect 56894 800 57002 856
rect 57170 800 57278 856
rect 57446 800 57554 856
rect 57722 800 57830 856
rect 57998 800 58106 856
rect 58274 800 58382 856
rect 58550 800 58658 856
rect 58826 800 58934 856
rect 59102 800 59210 856
rect 59378 800 59486 856
rect 59654 800 59762 856
rect 59930 800 60038 856
rect 60206 800 60314 856
rect 60482 800 60590 856
rect 60758 800 60866 856
rect 61034 800 61142 856
rect 61310 800 61418 856
rect 61586 800 61694 856
rect 61862 800 61970 856
rect 62138 800 62246 856
rect 62414 800 62522 856
rect 62690 800 62798 856
rect 62966 800 63074 856
rect 63242 800 63350 856
rect 63518 800 63626 856
rect 63794 800 63902 856
rect 64070 800 64178 856
rect 64346 800 64454 856
rect 64622 800 64730 856
rect 64898 800 65006 856
rect 65174 800 65282 856
rect 65450 800 65558 856
rect 65726 800 65834 856
rect 66002 800 66110 856
rect 66278 800 66386 856
rect 66554 800 66662 856
rect 66830 800 66938 856
rect 67106 800 67214 856
rect 67382 800 67490 856
rect 67658 800 67766 856
rect 67934 800 68042 856
rect 68210 800 68318 856
rect 68486 800 68594 856
rect 68762 800 68870 856
rect 69038 800 69146 856
rect 69314 800 69422 856
rect 69590 800 69698 856
rect 69866 800 69974 856
rect 70142 800 70250 856
rect 70418 800 70526 856
rect 70694 800 70802 856
rect 70970 800 71078 856
rect 71246 800 71354 856
rect 71522 800 71630 856
rect 71798 800 71906 856
rect 72074 800 72182 856
rect 72350 800 72458 856
rect 72626 800 72734 856
rect 72902 800 73010 856
rect 73178 800 73286 856
rect 73454 800 73562 856
rect 73730 800 73838 856
rect 74006 800 74114 856
rect 74282 800 74390 856
rect 74558 800 74666 856
rect 74834 800 74942 856
rect 75110 800 75218 856
rect 75386 800 75494 856
rect 75662 800 75770 856
rect 75938 800 76046 856
rect 76214 800 76322 856
rect 76490 800 76598 856
rect 76766 800 76874 856
rect 77042 800 77150 856
rect 77318 800 77426 856
rect 77594 800 77702 856
rect 77870 800 77978 856
rect 78146 800 78254 856
rect 78422 800 78530 856
rect 78698 800 78806 856
rect 78974 800 79082 856
rect 79250 800 79358 856
rect 79526 800 79634 856
rect 79802 800 79910 856
rect 80078 800 80186 856
rect 80354 800 80462 856
rect 80630 800 80738 856
rect 80906 800 81014 856
rect 81182 800 81290 856
rect 81458 800 81566 856
rect 81734 800 81842 856
rect 82010 800 82118 856
rect 82286 800 82394 856
rect 82562 800 82670 856
rect 82838 800 82946 856
rect 83114 800 83222 856
rect 83390 800 83498 856
rect 83666 800 83774 856
rect 83942 800 84050 856
rect 84218 800 84326 856
rect 84494 800 84602 856
rect 84770 800 84878 856
rect 85046 800 85154 856
rect 85322 800 85430 856
rect 85598 800 85706 856
rect 85874 800 85982 856
rect 86150 800 86258 856
rect 86426 800 86534 856
rect 86702 800 86810 856
rect 86978 800 87086 856
rect 87254 800 87362 856
rect 87530 800 87638 856
rect 87806 800 87914 856
rect 88082 800 88190 856
rect 88358 800 88466 856
rect 88634 800 88742 856
rect 88910 800 89018 856
rect 89186 800 89294 856
rect 89462 800 89570 856
rect 89738 800 89846 856
rect 90014 800 90122 856
rect 90290 800 90398 856
rect 90566 800 90674 856
rect 90842 800 90950 856
rect 91118 800 91226 856
rect 91394 800 91502 856
rect 91670 800 91778 856
rect 91946 800 92054 856
rect 92222 800 92330 856
rect 92498 800 92606 856
rect 92774 800 92882 856
rect 93050 800 93158 856
rect 93326 800 93434 856
rect 93602 800 93710 856
rect 93878 800 93986 856
rect 94154 800 94262 856
rect 94430 800 94538 856
rect 94706 800 94814 856
rect 94982 800 95090 856
rect 95258 800 95366 856
rect 95534 800 95642 856
rect 95810 800 95918 856
rect 96086 800 96194 856
rect 96362 800 96470 856
rect 96638 800 96746 856
rect 96914 800 97022 856
rect 97190 800 97298 856
rect 97466 800 97574 856
rect 97742 800 97850 856
rect 98018 800 98126 856
rect 98294 800 98402 856
rect 98570 800 98678 856
rect 98846 800 98954 856
rect 99122 800 99230 856
rect 99398 800 99506 856
rect 99674 800 99782 856
rect 99950 800 100058 856
rect 100226 800 100334 856
rect 100502 800 100610 856
rect 100778 800 100886 856
rect 101054 800 101162 856
rect 101330 800 101438 856
rect 101606 800 101714 856
rect 101882 800 101990 856
rect 102158 800 102266 856
rect 102434 800 102542 856
rect 102710 800 102818 856
rect 102986 800 103094 856
rect 103262 800 103370 856
rect 103538 800 103646 856
rect 103814 800 103922 856
rect 104090 800 104198 856
rect 104366 800 104474 856
rect 104642 800 104750 856
rect 104918 800 105026 856
rect 105194 800 105302 856
rect 105470 800 105578 856
rect 105746 800 105854 856
rect 106022 800 106130 856
rect 106298 800 106406 856
rect 106574 800 106682 856
rect 106850 800 106958 856
rect 107126 800 107234 856
rect 107402 800 107510 856
rect 107678 800 107786 856
rect 107954 800 108062 856
rect 108230 800 108338 856
rect 108506 800 108614 856
rect 108782 800 108890 856
rect 109058 800 109166 856
rect 109334 800 109442 856
rect 109610 800 109718 856
rect 109886 800 109994 856
rect 110162 800 110270 856
rect 110438 800 110546 856
rect 110714 800 110822 856
rect 110990 800 111098 856
rect 111266 800 111374 856
rect 111542 800 111650 856
rect 111818 800 111926 856
rect 112094 800 112202 856
rect 112370 800 112478 856
rect 112646 800 112754 856
rect 112922 800 113030 856
rect 113198 800 113306 856
rect 113474 800 113582 856
rect 113750 800 113858 856
rect 114026 800 114134 856
rect 114302 800 114410 856
rect 114578 800 114686 856
rect 114854 800 114962 856
rect 115130 800 115238 856
rect 115406 800 115514 856
rect 115682 800 115790 856
rect 115958 800 116066 856
rect 116234 800 116342 856
rect 116510 800 116618 856
rect 116786 800 116894 856
rect 117062 800 117170 856
rect 117338 800 117446 856
rect 117614 800 117722 856
rect 117890 800 117998 856
rect 118166 800 118274 856
rect 118442 800 118550 856
rect 118718 800 118826 856
rect 118994 800 119102 856
rect 119270 800 119378 856
rect 119546 800 119654 856
rect 119822 800 119930 856
rect 120098 800 120206 856
rect 120374 800 120482 856
rect 120650 800 120758 856
rect 120926 800 121034 856
rect 121202 800 121310 856
rect 121478 800 121586 856
rect 121754 800 121862 856
rect 122030 800 122138 856
rect 122306 800 122414 856
rect 122582 800 122690 856
rect 122858 800 122966 856
rect 123134 800 123242 856
rect 123410 800 123518 856
rect 123686 800 123794 856
rect 123962 800 124070 856
rect 124238 800 124346 856
rect 124514 800 124622 856
rect 124790 800 124898 856
rect 125066 800 125174 856
rect 125342 800 125450 856
rect 125618 800 125726 856
rect 125894 800 126002 856
rect 126170 800 126278 856
rect 126446 800 126554 856
rect 126722 800 126830 856
rect 126998 800 127106 856
rect 127274 800 127382 856
rect 127550 800 127658 856
rect 127826 800 127934 856
rect 128102 800 128210 856
rect 128378 800 128486 856
rect 128654 800 128762 856
rect 128930 800 129038 856
rect 129206 800 129314 856
rect 129482 800 129590 856
rect 129758 800 129866 856
rect 130034 800 130142 856
rect 130310 800 130418 856
rect 130586 800 130694 856
rect 130862 800 130970 856
rect 131138 800 131246 856
rect 131414 800 131522 856
rect 131690 800 131798 856
rect 131966 800 132074 856
rect 132242 800 132350 856
rect 132518 800 132626 856
rect 132794 800 132902 856
rect 133070 800 133178 856
rect 133346 800 133454 856
rect 133622 800 133730 856
rect 133898 800 134006 856
rect 134174 800 134282 856
rect 134450 800 134558 856
rect 134726 800 134834 856
rect 135002 800 135110 856
rect 135278 800 135386 856
rect 135554 800 135662 856
rect 135830 800 135938 856
<< metal3 >>
rect 135526 132200 136326 132320
rect 0 130024 800 130144
rect 0 127848 800 127968
rect 135526 127848 136326 127968
rect 0 125672 800 125792
rect 0 123496 800 123616
rect 135526 123496 136326 123616
rect 0 121320 800 121440
rect 0 119144 800 119264
rect 135526 119144 136326 119264
rect 0 116968 800 117088
rect 0 114792 800 114912
rect 135526 114792 136326 114912
rect 0 112616 800 112736
rect 0 110440 800 110560
rect 135526 110440 136326 110560
rect 0 108264 800 108384
rect 0 106088 800 106208
rect 135526 106088 136326 106208
rect 0 103912 800 104032
rect 0 101736 800 101856
rect 135526 101736 136326 101856
rect 0 99560 800 99680
rect 0 97384 800 97504
rect 135526 97384 136326 97504
rect 0 95208 800 95328
rect 0 93032 800 93152
rect 135526 93032 136326 93152
rect 0 90856 800 90976
rect 0 88680 800 88800
rect 135526 88680 136326 88800
rect 0 86504 800 86624
rect 0 84328 800 84448
rect 135526 84328 136326 84448
rect 0 82152 800 82272
rect 0 79976 800 80096
rect 135526 79976 136326 80096
rect 0 77800 800 77920
rect 0 75624 800 75744
rect 135526 75624 136326 75744
rect 0 73448 800 73568
rect 0 71272 800 71392
rect 135526 71272 136326 71392
rect 0 69096 800 69216
rect 0 66920 800 67040
rect 135526 66920 136326 67040
rect 0 64744 800 64864
rect 0 62568 800 62688
rect 135526 62568 136326 62688
rect 0 60392 800 60512
rect 0 58216 800 58336
rect 135526 58216 136326 58336
rect 0 56040 800 56160
rect 0 53864 800 53984
rect 135526 53864 136326 53984
rect 0 51688 800 51808
rect 0 49512 800 49632
rect 135526 49512 136326 49632
rect 0 47336 800 47456
rect 0 45160 800 45280
rect 135526 45160 136326 45280
rect 0 42984 800 43104
rect 0 40808 800 40928
rect 135526 40808 136326 40928
rect 0 38632 800 38752
rect 0 36456 800 36576
rect 135526 36456 136326 36576
rect 0 34280 800 34400
rect 0 32104 800 32224
rect 135526 32104 136326 32224
rect 0 29928 800 30048
rect 0 27752 800 27872
rect 135526 27752 136326 27872
rect 0 25576 800 25696
rect 0 23400 800 23520
rect 135526 23400 136326 23520
rect 0 21224 800 21344
rect 0 19048 800 19168
rect 135526 19048 136326 19168
rect 0 16872 800 16992
rect 0 14696 800 14816
rect 135526 14696 136326 14816
rect 0 12520 800 12640
rect 0 10344 800 10464
rect 135526 10344 136326 10464
rect 0 8168 800 8288
rect 135526 5992 136326 6112
<< obsm3 >>
rect 798 132400 135595 136033
rect 798 132120 135446 132400
rect 798 130224 135595 132120
rect 880 129944 135595 130224
rect 798 128048 135595 129944
rect 880 127768 135446 128048
rect 798 125872 135595 127768
rect 880 125592 135595 125872
rect 798 123696 135595 125592
rect 880 123416 135446 123696
rect 798 121520 135595 123416
rect 880 121240 135595 121520
rect 798 119344 135595 121240
rect 880 119064 135446 119344
rect 798 117168 135595 119064
rect 880 116888 135595 117168
rect 798 114992 135595 116888
rect 880 114712 135446 114992
rect 798 112816 135595 114712
rect 880 112536 135595 112816
rect 798 110640 135595 112536
rect 880 110360 135446 110640
rect 798 108464 135595 110360
rect 880 108184 135595 108464
rect 798 106288 135595 108184
rect 880 106008 135446 106288
rect 798 104112 135595 106008
rect 880 103832 135595 104112
rect 798 101936 135595 103832
rect 880 101656 135446 101936
rect 798 99760 135595 101656
rect 880 99480 135595 99760
rect 798 97584 135595 99480
rect 880 97304 135446 97584
rect 798 95408 135595 97304
rect 880 95128 135595 95408
rect 798 93232 135595 95128
rect 880 92952 135446 93232
rect 798 91056 135595 92952
rect 880 90776 135595 91056
rect 798 88880 135595 90776
rect 880 88600 135446 88880
rect 798 86704 135595 88600
rect 880 86424 135595 86704
rect 798 84528 135595 86424
rect 880 84248 135446 84528
rect 798 82352 135595 84248
rect 880 82072 135595 82352
rect 798 80176 135595 82072
rect 880 79896 135446 80176
rect 798 78000 135595 79896
rect 880 77720 135595 78000
rect 798 75824 135595 77720
rect 880 75544 135446 75824
rect 798 73648 135595 75544
rect 880 73368 135595 73648
rect 798 71472 135595 73368
rect 880 71192 135446 71472
rect 798 69296 135595 71192
rect 880 69016 135595 69296
rect 798 67120 135595 69016
rect 880 66840 135446 67120
rect 798 64944 135595 66840
rect 880 64664 135595 64944
rect 798 62768 135595 64664
rect 880 62488 135446 62768
rect 798 60592 135595 62488
rect 880 60312 135595 60592
rect 798 58416 135595 60312
rect 880 58136 135446 58416
rect 798 56240 135595 58136
rect 880 55960 135595 56240
rect 798 54064 135595 55960
rect 880 53784 135446 54064
rect 798 51888 135595 53784
rect 880 51608 135595 51888
rect 798 49712 135595 51608
rect 880 49432 135446 49712
rect 798 47536 135595 49432
rect 880 47256 135595 47536
rect 798 45360 135595 47256
rect 880 45080 135446 45360
rect 798 43184 135595 45080
rect 880 42904 135595 43184
rect 798 41008 135595 42904
rect 880 40728 135446 41008
rect 798 38832 135595 40728
rect 880 38552 135595 38832
rect 798 36656 135595 38552
rect 880 36376 135446 36656
rect 798 34480 135595 36376
rect 880 34200 135595 34480
rect 798 32304 135595 34200
rect 880 32024 135446 32304
rect 798 30128 135595 32024
rect 880 29848 135595 30128
rect 798 27952 135595 29848
rect 880 27672 135446 27952
rect 798 25776 135595 27672
rect 880 25496 135595 25776
rect 798 23600 135595 25496
rect 880 23320 135446 23600
rect 798 21424 135595 23320
rect 880 21144 135595 21424
rect 798 19248 135595 21144
rect 880 18968 135446 19248
rect 798 17072 135595 18968
rect 880 16792 135595 17072
rect 798 14896 135595 16792
rect 880 14616 135446 14896
rect 798 12720 135595 14616
rect 880 12440 135595 12720
rect 798 10544 135595 12440
rect 880 10264 135446 10544
rect 798 8368 135595 10264
rect 880 8088 135595 8368
rect 798 6192 135595 8088
rect 798 5912 135446 6192
rect 798 2143 135595 5912
<< metal4 >>
rect 3748 2128 4988 136048
rect 13748 2128 14988 136048
rect 23748 2128 24988 136048
rect 33748 2128 34988 136048
rect 43748 2128 44988 136048
rect 53748 2128 54988 136048
rect 63748 2128 64988 136048
rect 73748 2128 74988 136048
rect 83748 2128 84988 136048
rect 93748 2128 94988 136048
rect 103748 2128 104988 136048
rect 113748 2128 114988 136048
rect 123748 2128 124988 136048
rect 133748 2128 134988 136048
<< obsm4 >>
rect 10731 2347 13668 135285
rect 15068 2347 23668 135285
rect 25068 2347 33668 135285
rect 35068 2347 43668 135285
rect 45068 2347 53668 135285
rect 55068 2347 63668 135285
rect 65068 2347 73668 135285
rect 75068 2347 83668 135285
rect 85068 2347 93668 135285
rect 95068 2347 103668 135285
rect 105068 2347 113668 135285
rect 115068 2347 123668 135285
rect 125068 2347 133525 135285
<< labels >>
rlabel metal3 s 135526 5992 136326 6112 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 132682 137670 132738 138470 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 117778 137670 117834 138470 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 102874 137670 102930 138470 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 87970 137670 88026 138470 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 73066 137670 73122 138470 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 58162 137670 58218 138470 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 43258 137670 43314 138470 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 28354 137670 28410 138470 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 13450 137670 13506 138470 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 135526 19048 136326 19168 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 123496 800 123616 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 135526 32104 136326 32224 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 135526 45160 136326 45280 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 135526 58216 136326 58336 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 135526 71272 136326 71392 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 135526 84328 136326 84448 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 135526 97384 136326 97504 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 135526 110440 136326 110560 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 135526 123496 136326 123616 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 135526 14696 136326 14816 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 122746 137670 122802 138470 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 107842 137670 107898 138470 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 92938 137670 92994 138470 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 78034 137670 78090 138470 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 63130 137670 63186 138470 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 48226 137670 48282 138470 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 33322 137670 33378 138470 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 18418 137670 18474 138470 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 3514 137670 3570 138470 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 135526 27752 136326 27872 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 0 99560 800 99680 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 93032 800 93152 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 86504 800 86624 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 66920 800 67040 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 135526 40808 136326 40928 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 135526 53864 136326 53984 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 135526 66920 136326 67040 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 135526 79976 136326 80096 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 135526 93032 136326 93152 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 135526 106088 136326 106208 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 135526 119144 136326 119264 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 135526 132200 136326 132320 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 135526 10344 136326 10464 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 127714 137670 127770 138470 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 112810 137670 112866 138470 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 97906 137670 97962 138470 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 83002 137670 83058 138470 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 68098 137670 68154 138470 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 53194 137670 53250 138470 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 38290 137670 38346 138470 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 23386 137670 23442 138470 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 8482 137670 8538 138470 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 135526 23400 136326 23520 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 0 121320 800 121440 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 0 108264 800 108384 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 0 101736 800 101856 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 88680 800 88800 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 82152 800 82272 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 69096 800 69216 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 135526 36456 136326 36576 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 135526 49512 136326 49632 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 135526 62568 136326 62688 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 135526 75624 136326 75744 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 135526 88680 136326 88800 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 135526 101736 136326 101856 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 135526 114792 136326 114912 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 135526 127848 136326 127968 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 133234 0 133290 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 134890 0 134946 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 3748 2128 4988 136048 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 23748 2128 24988 136048 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 43748 2128 44988 136048 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 63748 2128 64988 136048 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 83748 2128 84988 136048 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 103748 2128 104988 136048 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 123748 2128 124988 136048 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 13748 2128 14988 136048 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 33748 2128 34988 136048 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 53748 2128 54988 136048 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 73748 2128 74988 136048 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 93748 2128 94988 136048 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 113748 2128 114988 136048 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 133748 2128 134988 136048 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 478 0 534 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 136326 138470
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 68997724
string GDS_FILE /home/ejjimenezu/Repos/caravel_simple_fpu/openlane/fpu/runs/24_12_05_02_02/results/signoff/fpu.magic.gds
string GDS_START 1076512
<< end >>

