magic
tech sky130A
magscale 1 2
timestamp 1733317639
<< obsli1 >>
rect 1104 2159 142600 143633
<< obsm1 >>
rect 934 1232 142660 143664
<< metal2 >>
rect 3698 145109 3754 145909
rect 8942 145109 8998 145909
rect 14186 145109 14242 145909
rect 19430 145109 19486 145909
rect 24674 145109 24730 145909
rect 29918 145109 29974 145909
rect 35162 145109 35218 145909
rect 40406 145109 40462 145909
rect 45650 145109 45706 145909
rect 50894 145109 50950 145909
rect 56138 145109 56194 145909
rect 61382 145109 61438 145909
rect 66626 145109 66682 145909
rect 71870 145109 71926 145909
rect 77114 145109 77170 145909
rect 82358 145109 82414 145909
rect 87602 145109 87658 145909
rect 92846 145109 92902 145909
rect 98090 145109 98146 145909
rect 103334 145109 103390 145909
rect 108578 145109 108634 145909
rect 113822 145109 113878 145909
rect 119066 145109 119122 145909
rect 124310 145109 124366 145909
rect 129554 145109 129610 145909
rect 134798 145109 134854 145909
rect 140042 145109 140098 145909
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54758 0 54814 800
rect 55034 0 55090 800
rect 55310 0 55366 800
rect 55586 0 55642 800
rect 55862 0 55918 800
rect 56138 0 56194 800
rect 56414 0 56470 800
rect 56690 0 56746 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58622 0 58678 800
rect 58898 0 58954 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59726 0 59782 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61382 0 61438 800
rect 61658 0 61714 800
rect 61934 0 61990 800
rect 62210 0 62266 800
rect 62486 0 62542 800
rect 62762 0 62818 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63590 0 63646 800
rect 63866 0 63922 800
rect 64142 0 64198 800
rect 64418 0 64474 800
rect 64694 0 64750 800
rect 64970 0 65026 800
rect 65246 0 65302 800
rect 65522 0 65578 800
rect 65798 0 65854 800
rect 66074 0 66130 800
rect 66350 0 66406 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 68006 0 68062 800
rect 68282 0 68338 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69110 0 69166 800
rect 69386 0 69442 800
rect 69662 0 69718 800
rect 69938 0 69994 800
rect 70214 0 70270 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 71042 0 71098 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71870 0 71926 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72698 0 72754 800
rect 72974 0 73030 800
rect 73250 0 73306 800
rect 73526 0 73582 800
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75182 0 75238 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 76010 0 76066 800
rect 76286 0 76342 800
rect 76562 0 76618 800
rect 76838 0 76894 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78770 0 78826 800
rect 79046 0 79102 800
rect 79322 0 79378 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80150 0 80206 800
rect 80426 0 80482 800
rect 80702 0 80758 800
rect 80978 0 81034 800
rect 81254 0 81310 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 82082 0 82138 800
rect 82358 0 82414 800
rect 82634 0 82690 800
rect 82910 0 82966 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83738 0 83794 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84566 0 84622 800
rect 84842 0 84898 800
rect 85118 0 85174 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 85946 0 86002 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86774 0 86830 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87602 0 87658 800
rect 87878 0 87934 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88706 0 88762 800
rect 88982 0 89038 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89810 0 89866 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90638 0 90694 800
rect 90914 0 90970 800
rect 91190 0 91246 800
rect 91466 0 91522 800
rect 91742 0 91798 800
rect 92018 0 92074 800
rect 92294 0 92350 800
rect 92570 0 92626 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93674 0 93730 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94502 0 94558 800
rect 94778 0 94834 800
rect 95054 0 95110 800
rect 95330 0 95386 800
rect 95606 0 95662 800
rect 95882 0 95938 800
rect 96158 0 96214 800
rect 96434 0 96490 800
rect 96710 0 96766 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97538 0 97594 800
rect 97814 0 97870 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99194 0 99250 800
rect 99470 0 99526 800
rect 99746 0 99802 800
rect 100022 0 100078 800
rect 100298 0 100354 800
rect 100574 0 100630 800
rect 100850 0 100906 800
rect 101126 0 101182 800
rect 101402 0 101458 800
rect 101678 0 101734 800
rect 101954 0 102010 800
rect 102230 0 102286 800
rect 102506 0 102562 800
rect 102782 0 102838 800
rect 103058 0 103114 800
rect 103334 0 103390 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104714 0 104770 800
rect 104990 0 105046 800
rect 105266 0 105322 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106094 0 106150 800
rect 106370 0 106426 800
rect 106646 0 106702 800
rect 106922 0 106978 800
rect 107198 0 107254 800
rect 107474 0 107530 800
rect 107750 0 107806 800
rect 108026 0 108082 800
rect 108302 0 108358 800
rect 108578 0 108634 800
rect 108854 0 108910 800
rect 109130 0 109186 800
rect 109406 0 109462 800
rect 109682 0 109738 800
rect 109958 0 110014 800
rect 110234 0 110290 800
rect 110510 0 110566 800
rect 110786 0 110842 800
rect 111062 0 111118 800
rect 111338 0 111394 800
rect 111614 0 111670 800
rect 111890 0 111946 800
rect 112166 0 112222 800
rect 112442 0 112498 800
rect 112718 0 112774 800
rect 112994 0 113050 800
rect 113270 0 113326 800
rect 113546 0 113602 800
rect 113822 0 113878 800
rect 114098 0 114154 800
rect 114374 0 114430 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115202 0 115258 800
rect 115478 0 115534 800
rect 115754 0 115810 800
rect 116030 0 116086 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117134 0 117190 800
rect 117410 0 117466 800
rect 117686 0 117742 800
rect 117962 0 118018 800
rect 118238 0 118294 800
rect 118514 0 118570 800
rect 118790 0 118846 800
rect 119066 0 119122 800
rect 119342 0 119398 800
rect 119618 0 119674 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120446 0 120502 800
rect 120722 0 120778 800
rect 120998 0 121054 800
rect 121274 0 121330 800
rect 121550 0 121606 800
rect 121826 0 121882 800
rect 122102 0 122158 800
rect 122378 0 122434 800
rect 122654 0 122710 800
rect 122930 0 122986 800
rect 123206 0 123262 800
rect 123482 0 123538 800
rect 123758 0 123814 800
rect 124034 0 124090 800
rect 124310 0 124366 800
rect 124586 0 124642 800
rect 124862 0 124918 800
rect 125138 0 125194 800
rect 125414 0 125470 800
rect 125690 0 125746 800
rect 125966 0 126022 800
rect 126242 0 126298 800
rect 126518 0 126574 800
rect 126794 0 126850 800
rect 127070 0 127126 800
rect 127346 0 127402 800
rect 127622 0 127678 800
rect 127898 0 127954 800
rect 128174 0 128230 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129002 0 129058 800
rect 129278 0 129334 800
rect 129554 0 129610 800
rect 129830 0 129886 800
rect 130106 0 130162 800
rect 130382 0 130438 800
rect 130658 0 130714 800
rect 130934 0 130990 800
rect 131210 0 131266 800
rect 131486 0 131542 800
rect 131762 0 131818 800
rect 132038 0 132094 800
rect 132314 0 132370 800
rect 132590 0 132646 800
rect 132866 0 132922 800
rect 133142 0 133198 800
rect 133418 0 133474 800
rect 133694 0 133750 800
rect 133970 0 134026 800
rect 134246 0 134302 800
rect 134522 0 134578 800
rect 134798 0 134854 800
rect 135074 0 135130 800
rect 135350 0 135406 800
rect 135626 0 135682 800
rect 135902 0 135958 800
rect 136178 0 136234 800
rect 136454 0 136510 800
rect 136730 0 136786 800
rect 137006 0 137062 800
rect 137282 0 137338 800
rect 137558 0 137614 800
rect 137834 0 137890 800
rect 138110 0 138166 800
rect 138386 0 138442 800
rect 138662 0 138718 800
rect 138938 0 138994 800
rect 139214 0 139270 800
rect 139490 0 139546 800
rect 139766 0 139822 800
<< obsm2 >>
rect 938 145053 3642 145194
rect 3810 145053 8886 145194
rect 9054 145053 14130 145194
rect 14298 145053 19374 145194
rect 19542 145053 24618 145194
rect 24786 145053 29862 145194
rect 30030 145053 35106 145194
rect 35274 145053 40350 145194
rect 40518 145053 45594 145194
rect 45762 145053 50838 145194
rect 51006 145053 56082 145194
rect 56250 145053 61326 145194
rect 61494 145053 66570 145194
rect 66738 145053 71814 145194
rect 71982 145053 77058 145194
rect 77226 145053 82302 145194
rect 82470 145053 87546 145194
rect 87714 145053 92790 145194
rect 92958 145053 98034 145194
rect 98202 145053 103278 145194
rect 103446 145053 108522 145194
rect 108690 145053 113766 145194
rect 113934 145053 119010 145194
rect 119178 145053 124254 145194
rect 124422 145053 129498 145194
rect 129666 145053 134742 145194
rect 134910 145053 139986 145194
rect 140154 145053 142582 145194
rect 938 856 142582 145053
rect 938 734 3918 856
rect 4086 734 4194 856
rect 4362 734 4470 856
rect 4638 734 4746 856
rect 4914 734 5022 856
rect 5190 734 5298 856
rect 5466 734 5574 856
rect 5742 734 5850 856
rect 6018 734 6126 856
rect 6294 734 6402 856
rect 6570 734 6678 856
rect 6846 734 6954 856
rect 7122 734 7230 856
rect 7398 734 7506 856
rect 7674 734 7782 856
rect 7950 734 8058 856
rect 8226 734 8334 856
rect 8502 734 8610 856
rect 8778 734 8886 856
rect 9054 734 9162 856
rect 9330 734 9438 856
rect 9606 734 9714 856
rect 9882 734 9990 856
rect 10158 734 10266 856
rect 10434 734 10542 856
rect 10710 734 10818 856
rect 10986 734 11094 856
rect 11262 734 11370 856
rect 11538 734 11646 856
rect 11814 734 11922 856
rect 12090 734 12198 856
rect 12366 734 12474 856
rect 12642 734 12750 856
rect 12918 734 13026 856
rect 13194 734 13302 856
rect 13470 734 13578 856
rect 13746 734 13854 856
rect 14022 734 14130 856
rect 14298 734 14406 856
rect 14574 734 14682 856
rect 14850 734 14958 856
rect 15126 734 15234 856
rect 15402 734 15510 856
rect 15678 734 15786 856
rect 15954 734 16062 856
rect 16230 734 16338 856
rect 16506 734 16614 856
rect 16782 734 16890 856
rect 17058 734 17166 856
rect 17334 734 17442 856
rect 17610 734 17718 856
rect 17886 734 17994 856
rect 18162 734 18270 856
rect 18438 734 18546 856
rect 18714 734 18822 856
rect 18990 734 19098 856
rect 19266 734 19374 856
rect 19542 734 19650 856
rect 19818 734 19926 856
rect 20094 734 20202 856
rect 20370 734 20478 856
rect 20646 734 20754 856
rect 20922 734 21030 856
rect 21198 734 21306 856
rect 21474 734 21582 856
rect 21750 734 21858 856
rect 22026 734 22134 856
rect 22302 734 22410 856
rect 22578 734 22686 856
rect 22854 734 22962 856
rect 23130 734 23238 856
rect 23406 734 23514 856
rect 23682 734 23790 856
rect 23958 734 24066 856
rect 24234 734 24342 856
rect 24510 734 24618 856
rect 24786 734 24894 856
rect 25062 734 25170 856
rect 25338 734 25446 856
rect 25614 734 25722 856
rect 25890 734 25998 856
rect 26166 734 26274 856
rect 26442 734 26550 856
rect 26718 734 26826 856
rect 26994 734 27102 856
rect 27270 734 27378 856
rect 27546 734 27654 856
rect 27822 734 27930 856
rect 28098 734 28206 856
rect 28374 734 28482 856
rect 28650 734 28758 856
rect 28926 734 29034 856
rect 29202 734 29310 856
rect 29478 734 29586 856
rect 29754 734 29862 856
rect 30030 734 30138 856
rect 30306 734 30414 856
rect 30582 734 30690 856
rect 30858 734 30966 856
rect 31134 734 31242 856
rect 31410 734 31518 856
rect 31686 734 31794 856
rect 31962 734 32070 856
rect 32238 734 32346 856
rect 32514 734 32622 856
rect 32790 734 32898 856
rect 33066 734 33174 856
rect 33342 734 33450 856
rect 33618 734 33726 856
rect 33894 734 34002 856
rect 34170 734 34278 856
rect 34446 734 34554 856
rect 34722 734 34830 856
rect 34998 734 35106 856
rect 35274 734 35382 856
rect 35550 734 35658 856
rect 35826 734 35934 856
rect 36102 734 36210 856
rect 36378 734 36486 856
rect 36654 734 36762 856
rect 36930 734 37038 856
rect 37206 734 37314 856
rect 37482 734 37590 856
rect 37758 734 37866 856
rect 38034 734 38142 856
rect 38310 734 38418 856
rect 38586 734 38694 856
rect 38862 734 38970 856
rect 39138 734 39246 856
rect 39414 734 39522 856
rect 39690 734 39798 856
rect 39966 734 40074 856
rect 40242 734 40350 856
rect 40518 734 40626 856
rect 40794 734 40902 856
rect 41070 734 41178 856
rect 41346 734 41454 856
rect 41622 734 41730 856
rect 41898 734 42006 856
rect 42174 734 42282 856
rect 42450 734 42558 856
rect 42726 734 42834 856
rect 43002 734 43110 856
rect 43278 734 43386 856
rect 43554 734 43662 856
rect 43830 734 43938 856
rect 44106 734 44214 856
rect 44382 734 44490 856
rect 44658 734 44766 856
rect 44934 734 45042 856
rect 45210 734 45318 856
rect 45486 734 45594 856
rect 45762 734 45870 856
rect 46038 734 46146 856
rect 46314 734 46422 856
rect 46590 734 46698 856
rect 46866 734 46974 856
rect 47142 734 47250 856
rect 47418 734 47526 856
rect 47694 734 47802 856
rect 47970 734 48078 856
rect 48246 734 48354 856
rect 48522 734 48630 856
rect 48798 734 48906 856
rect 49074 734 49182 856
rect 49350 734 49458 856
rect 49626 734 49734 856
rect 49902 734 50010 856
rect 50178 734 50286 856
rect 50454 734 50562 856
rect 50730 734 50838 856
rect 51006 734 51114 856
rect 51282 734 51390 856
rect 51558 734 51666 856
rect 51834 734 51942 856
rect 52110 734 52218 856
rect 52386 734 52494 856
rect 52662 734 52770 856
rect 52938 734 53046 856
rect 53214 734 53322 856
rect 53490 734 53598 856
rect 53766 734 53874 856
rect 54042 734 54150 856
rect 54318 734 54426 856
rect 54594 734 54702 856
rect 54870 734 54978 856
rect 55146 734 55254 856
rect 55422 734 55530 856
rect 55698 734 55806 856
rect 55974 734 56082 856
rect 56250 734 56358 856
rect 56526 734 56634 856
rect 56802 734 56910 856
rect 57078 734 57186 856
rect 57354 734 57462 856
rect 57630 734 57738 856
rect 57906 734 58014 856
rect 58182 734 58290 856
rect 58458 734 58566 856
rect 58734 734 58842 856
rect 59010 734 59118 856
rect 59286 734 59394 856
rect 59562 734 59670 856
rect 59838 734 59946 856
rect 60114 734 60222 856
rect 60390 734 60498 856
rect 60666 734 60774 856
rect 60942 734 61050 856
rect 61218 734 61326 856
rect 61494 734 61602 856
rect 61770 734 61878 856
rect 62046 734 62154 856
rect 62322 734 62430 856
rect 62598 734 62706 856
rect 62874 734 62982 856
rect 63150 734 63258 856
rect 63426 734 63534 856
rect 63702 734 63810 856
rect 63978 734 64086 856
rect 64254 734 64362 856
rect 64530 734 64638 856
rect 64806 734 64914 856
rect 65082 734 65190 856
rect 65358 734 65466 856
rect 65634 734 65742 856
rect 65910 734 66018 856
rect 66186 734 66294 856
rect 66462 734 66570 856
rect 66738 734 66846 856
rect 67014 734 67122 856
rect 67290 734 67398 856
rect 67566 734 67674 856
rect 67842 734 67950 856
rect 68118 734 68226 856
rect 68394 734 68502 856
rect 68670 734 68778 856
rect 68946 734 69054 856
rect 69222 734 69330 856
rect 69498 734 69606 856
rect 69774 734 69882 856
rect 70050 734 70158 856
rect 70326 734 70434 856
rect 70602 734 70710 856
rect 70878 734 70986 856
rect 71154 734 71262 856
rect 71430 734 71538 856
rect 71706 734 71814 856
rect 71982 734 72090 856
rect 72258 734 72366 856
rect 72534 734 72642 856
rect 72810 734 72918 856
rect 73086 734 73194 856
rect 73362 734 73470 856
rect 73638 734 73746 856
rect 73914 734 74022 856
rect 74190 734 74298 856
rect 74466 734 74574 856
rect 74742 734 74850 856
rect 75018 734 75126 856
rect 75294 734 75402 856
rect 75570 734 75678 856
rect 75846 734 75954 856
rect 76122 734 76230 856
rect 76398 734 76506 856
rect 76674 734 76782 856
rect 76950 734 77058 856
rect 77226 734 77334 856
rect 77502 734 77610 856
rect 77778 734 77886 856
rect 78054 734 78162 856
rect 78330 734 78438 856
rect 78606 734 78714 856
rect 78882 734 78990 856
rect 79158 734 79266 856
rect 79434 734 79542 856
rect 79710 734 79818 856
rect 79986 734 80094 856
rect 80262 734 80370 856
rect 80538 734 80646 856
rect 80814 734 80922 856
rect 81090 734 81198 856
rect 81366 734 81474 856
rect 81642 734 81750 856
rect 81918 734 82026 856
rect 82194 734 82302 856
rect 82470 734 82578 856
rect 82746 734 82854 856
rect 83022 734 83130 856
rect 83298 734 83406 856
rect 83574 734 83682 856
rect 83850 734 83958 856
rect 84126 734 84234 856
rect 84402 734 84510 856
rect 84678 734 84786 856
rect 84954 734 85062 856
rect 85230 734 85338 856
rect 85506 734 85614 856
rect 85782 734 85890 856
rect 86058 734 86166 856
rect 86334 734 86442 856
rect 86610 734 86718 856
rect 86886 734 86994 856
rect 87162 734 87270 856
rect 87438 734 87546 856
rect 87714 734 87822 856
rect 87990 734 88098 856
rect 88266 734 88374 856
rect 88542 734 88650 856
rect 88818 734 88926 856
rect 89094 734 89202 856
rect 89370 734 89478 856
rect 89646 734 89754 856
rect 89922 734 90030 856
rect 90198 734 90306 856
rect 90474 734 90582 856
rect 90750 734 90858 856
rect 91026 734 91134 856
rect 91302 734 91410 856
rect 91578 734 91686 856
rect 91854 734 91962 856
rect 92130 734 92238 856
rect 92406 734 92514 856
rect 92682 734 92790 856
rect 92958 734 93066 856
rect 93234 734 93342 856
rect 93510 734 93618 856
rect 93786 734 93894 856
rect 94062 734 94170 856
rect 94338 734 94446 856
rect 94614 734 94722 856
rect 94890 734 94998 856
rect 95166 734 95274 856
rect 95442 734 95550 856
rect 95718 734 95826 856
rect 95994 734 96102 856
rect 96270 734 96378 856
rect 96546 734 96654 856
rect 96822 734 96930 856
rect 97098 734 97206 856
rect 97374 734 97482 856
rect 97650 734 97758 856
rect 97926 734 98034 856
rect 98202 734 98310 856
rect 98478 734 98586 856
rect 98754 734 98862 856
rect 99030 734 99138 856
rect 99306 734 99414 856
rect 99582 734 99690 856
rect 99858 734 99966 856
rect 100134 734 100242 856
rect 100410 734 100518 856
rect 100686 734 100794 856
rect 100962 734 101070 856
rect 101238 734 101346 856
rect 101514 734 101622 856
rect 101790 734 101898 856
rect 102066 734 102174 856
rect 102342 734 102450 856
rect 102618 734 102726 856
rect 102894 734 103002 856
rect 103170 734 103278 856
rect 103446 734 103554 856
rect 103722 734 103830 856
rect 103998 734 104106 856
rect 104274 734 104382 856
rect 104550 734 104658 856
rect 104826 734 104934 856
rect 105102 734 105210 856
rect 105378 734 105486 856
rect 105654 734 105762 856
rect 105930 734 106038 856
rect 106206 734 106314 856
rect 106482 734 106590 856
rect 106758 734 106866 856
rect 107034 734 107142 856
rect 107310 734 107418 856
rect 107586 734 107694 856
rect 107862 734 107970 856
rect 108138 734 108246 856
rect 108414 734 108522 856
rect 108690 734 108798 856
rect 108966 734 109074 856
rect 109242 734 109350 856
rect 109518 734 109626 856
rect 109794 734 109902 856
rect 110070 734 110178 856
rect 110346 734 110454 856
rect 110622 734 110730 856
rect 110898 734 111006 856
rect 111174 734 111282 856
rect 111450 734 111558 856
rect 111726 734 111834 856
rect 112002 734 112110 856
rect 112278 734 112386 856
rect 112554 734 112662 856
rect 112830 734 112938 856
rect 113106 734 113214 856
rect 113382 734 113490 856
rect 113658 734 113766 856
rect 113934 734 114042 856
rect 114210 734 114318 856
rect 114486 734 114594 856
rect 114762 734 114870 856
rect 115038 734 115146 856
rect 115314 734 115422 856
rect 115590 734 115698 856
rect 115866 734 115974 856
rect 116142 734 116250 856
rect 116418 734 116526 856
rect 116694 734 116802 856
rect 116970 734 117078 856
rect 117246 734 117354 856
rect 117522 734 117630 856
rect 117798 734 117906 856
rect 118074 734 118182 856
rect 118350 734 118458 856
rect 118626 734 118734 856
rect 118902 734 119010 856
rect 119178 734 119286 856
rect 119454 734 119562 856
rect 119730 734 119838 856
rect 120006 734 120114 856
rect 120282 734 120390 856
rect 120558 734 120666 856
rect 120834 734 120942 856
rect 121110 734 121218 856
rect 121386 734 121494 856
rect 121662 734 121770 856
rect 121938 734 122046 856
rect 122214 734 122322 856
rect 122490 734 122598 856
rect 122766 734 122874 856
rect 123042 734 123150 856
rect 123318 734 123426 856
rect 123594 734 123702 856
rect 123870 734 123978 856
rect 124146 734 124254 856
rect 124422 734 124530 856
rect 124698 734 124806 856
rect 124974 734 125082 856
rect 125250 734 125358 856
rect 125526 734 125634 856
rect 125802 734 125910 856
rect 126078 734 126186 856
rect 126354 734 126462 856
rect 126630 734 126738 856
rect 126906 734 127014 856
rect 127182 734 127290 856
rect 127458 734 127566 856
rect 127734 734 127842 856
rect 128010 734 128118 856
rect 128286 734 128394 856
rect 128562 734 128670 856
rect 128838 734 128946 856
rect 129114 734 129222 856
rect 129390 734 129498 856
rect 129666 734 129774 856
rect 129942 734 130050 856
rect 130218 734 130326 856
rect 130494 734 130602 856
rect 130770 734 130878 856
rect 131046 734 131154 856
rect 131322 734 131430 856
rect 131598 734 131706 856
rect 131874 734 131982 856
rect 132150 734 132258 856
rect 132426 734 132534 856
rect 132702 734 132810 856
rect 132978 734 133086 856
rect 133254 734 133362 856
rect 133530 734 133638 856
rect 133806 734 133914 856
rect 134082 734 134190 856
rect 134358 734 134466 856
rect 134634 734 134742 856
rect 134910 734 135018 856
rect 135186 734 135294 856
rect 135462 734 135570 856
rect 135738 734 135846 856
rect 136014 734 136122 856
rect 136290 734 136398 856
rect 136566 734 136674 856
rect 136842 734 136950 856
rect 137118 734 137226 856
rect 137394 734 137502 856
rect 137670 734 137778 856
rect 137946 734 138054 856
rect 138222 734 138330 856
rect 138498 734 138606 856
rect 138774 734 138882 856
rect 139050 734 139158 856
rect 139326 734 139434 856
rect 139602 734 139710 856
rect 139878 734 142582 856
<< metal3 >>
rect 0 141448 800 141568
rect 142965 139816 143765 139936
rect 0 139000 800 139120
rect 0 136552 800 136672
rect 142965 135192 143765 135312
rect 0 134104 800 134224
rect 0 131656 800 131776
rect 142965 130568 143765 130688
rect 0 129208 800 129328
rect 0 126760 800 126880
rect 142965 125944 143765 126064
rect 0 124312 800 124432
rect 0 121864 800 121984
rect 142965 121320 143765 121440
rect 0 119416 800 119536
rect 0 116968 800 117088
rect 142965 116696 143765 116816
rect 0 114520 800 114640
rect 0 112072 800 112192
rect 142965 112072 143765 112192
rect 0 109624 800 109744
rect 142965 107448 143765 107568
rect 0 107176 800 107296
rect 0 104728 800 104848
rect 142965 102824 143765 102944
rect 0 102280 800 102400
rect 0 99832 800 99952
rect 142965 98200 143765 98320
rect 0 97384 800 97504
rect 0 94936 800 95056
rect 142965 93576 143765 93696
rect 0 92488 800 92608
rect 0 90040 800 90160
rect 142965 88952 143765 89072
rect 0 87592 800 87712
rect 0 85144 800 85264
rect 142965 84328 143765 84448
rect 0 82696 800 82816
rect 0 80248 800 80368
rect 142965 79704 143765 79824
rect 0 77800 800 77920
rect 0 75352 800 75472
rect 142965 75080 143765 75200
rect 0 72904 800 73024
rect 0 70456 800 70576
rect 142965 70456 143765 70576
rect 0 68008 800 68128
rect 142965 65832 143765 65952
rect 0 65560 800 65680
rect 0 63112 800 63232
rect 142965 61208 143765 61328
rect 0 60664 800 60784
rect 0 58216 800 58336
rect 142965 56584 143765 56704
rect 0 55768 800 55888
rect 0 53320 800 53440
rect 142965 51960 143765 52080
rect 0 50872 800 50992
rect 0 48424 800 48544
rect 142965 47336 143765 47456
rect 0 45976 800 46096
rect 0 43528 800 43648
rect 142965 42712 143765 42832
rect 0 41080 800 41200
rect 0 38632 800 38752
rect 142965 38088 143765 38208
rect 0 36184 800 36304
rect 0 33736 800 33856
rect 142965 33464 143765 33584
rect 0 31288 800 31408
rect 0 28840 800 28960
rect 142965 28840 143765 28960
rect 0 26392 800 26512
rect 142965 24216 143765 24336
rect 0 23944 800 24064
rect 0 21496 800 21616
rect 142965 19592 143765 19712
rect 0 19048 800 19168
rect 0 16600 800 16720
rect 142965 14968 143765 15088
rect 0 14152 800 14272
rect 0 11704 800 11824
rect 142965 10344 143765 10464
rect 0 9256 800 9376
rect 0 6808 800 6928
rect 142965 5720 143765 5840
rect 0 4360 800 4480
<< obsm3 >>
rect 798 141648 142965 143649
rect 880 141368 142965 141648
rect 798 140016 142965 141368
rect 798 139736 142885 140016
rect 798 139200 142965 139736
rect 880 138920 142965 139200
rect 798 136752 142965 138920
rect 880 136472 142965 136752
rect 798 135392 142965 136472
rect 798 135112 142885 135392
rect 798 134304 142965 135112
rect 880 134024 142965 134304
rect 798 131856 142965 134024
rect 880 131576 142965 131856
rect 798 130768 142965 131576
rect 798 130488 142885 130768
rect 798 129408 142965 130488
rect 880 129128 142965 129408
rect 798 126960 142965 129128
rect 880 126680 142965 126960
rect 798 126144 142965 126680
rect 798 125864 142885 126144
rect 798 124512 142965 125864
rect 880 124232 142965 124512
rect 798 122064 142965 124232
rect 880 121784 142965 122064
rect 798 121520 142965 121784
rect 798 121240 142885 121520
rect 798 119616 142965 121240
rect 880 119336 142965 119616
rect 798 117168 142965 119336
rect 880 116896 142965 117168
rect 880 116888 142885 116896
rect 798 116616 142885 116888
rect 798 114720 142965 116616
rect 880 114440 142965 114720
rect 798 112272 142965 114440
rect 880 111992 142885 112272
rect 798 109824 142965 111992
rect 880 109544 142965 109824
rect 798 107648 142965 109544
rect 798 107376 142885 107648
rect 880 107368 142885 107376
rect 880 107096 142965 107368
rect 798 104928 142965 107096
rect 880 104648 142965 104928
rect 798 103024 142965 104648
rect 798 102744 142885 103024
rect 798 102480 142965 102744
rect 880 102200 142965 102480
rect 798 100032 142965 102200
rect 880 99752 142965 100032
rect 798 98400 142965 99752
rect 798 98120 142885 98400
rect 798 97584 142965 98120
rect 880 97304 142965 97584
rect 798 95136 142965 97304
rect 880 94856 142965 95136
rect 798 93776 142965 94856
rect 798 93496 142885 93776
rect 798 92688 142965 93496
rect 880 92408 142965 92688
rect 798 90240 142965 92408
rect 880 89960 142965 90240
rect 798 89152 142965 89960
rect 798 88872 142885 89152
rect 798 87792 142965 88872
rect 880 87512 142965 87792
rect 798 85344 142965 87512
rect 880 85064 142965 85344
rect 798 84528 142965 85064
rect 798 84248 142885 84528
rect 798 82896 142965 84248
rect 880 82616 142965 82896
rect 798 80448 142965 82616
rect 880 80168 142965 80448
rect 798 79904 142965 80168
rect 798 79624 142885 79904
rect 798 78000 142965 79624
rect 880 77720 142965 78000
rect 798 75552 142965 77720
rect 880 75280 142965 75552
rect 880 75272 142885 75280
rect 798 75000 142885 75272
rect 798 73104 142965 75000
rect 880 72824 142965 73104
rect 798 70656 142965 72824
rect 880 70376 142885 70656
rect 798 68208 142965 70376
rect 880 67928 142965 68208
rect 798 66032 142965 67928
rect 798 65760 142885 66032
rect 880 65752 142885 65760
rect 880 65480 142965 65752
rect 798 63312 142965 65480
rect 880 63032 142965 63312
rect 798 61408 142965 63032
rect 798 61128 142885 61408
rect 798 60864 142965 61128
rect 880 60584 142965 60864
rect 798 58416 142965 60584
rect 880 58136 142965 58416
rect 798 56784 142965 58136
rect 798 56504 142885 56784
rect 798 55968 142965 56504
rect 880 55688 142965 55968
rect 798 53520 142965 55688
rect 880 53240 142965 53520
rect 798 52160 142965 53240
rect 798 51880 142885 52160
rect 798 51072 142965 51880
rect 880 50792 142965 51072
rect 798 48624 142965 50792
rect 880 48344 142965 48624
rect 798 47536 142965 48344
rect 798 47256 142885 47536
rect 798 46176 142965 47256
rect 880 45896 142965 46176
rect 798 43728 142965 45896
rect 880 43448 142965 43728
rect 798 42912 142965 43448
rect 798 42632 142885 42912
rect 798 41280 142965 42632
rect 880 41000 142965 41280
rect 798 38832 142965 41000
rect 880 38552 142965 38832
rect 798 38288 142965 38552
rect 798 38008 142885 38288
rect 798 36384 142965 38008
rect 880 36104 142965 36384
rect 798 33936 142965 36104
rect 880 33664 142965 33936
rect 880 33656 142885 33664
rect 798 33384 142885 33656
rect 798 31488 142965 33384
rect 880 31208 142965 31488
rect 798 29040 142965 31208
rect 880 28760 142885 29040
rect 798 26592 142965 28760
rect 880 26312 142965 26592
rect 798 24416 142965 26312
rect 798 24144 142885 24416
rect 880 24136 142885 24144
rect 880 23864 142965 24136
rect 798 21696 142965 23864
rect 880 21416 142965 21696
rect 798 19792 142965 21416
rect 798 19512 142885 19792
rect 798 19248 142965 19512
rect 880 18968 142965 19248
rect 798 16800 142965 18968
rect 880 16520 142965 16800
rect 798 15168 142965 16520
rect 798 14888 142885 15168
rect 798 14352 142965 14888
rect 880 14072 142965 14352
rect 798 11904 142965 14072
rect 880 11624 142965 11904
rect 798 10544 142965 11624
rect 798 10264 142885 10544
rect 798 9456 142965 10264
rect 880 9176 142965 9456
rect 798 7008 142965 9176
rect 880 6728 142965 7008
rect 798 5920 142965 6728
rect 798 5640 142885 5920
rect 798 4560 142965 5640
rect 880 4280 142965 4560
rect 798 2143 142965 4280
<< metal4 >>
rect 3748 2128 4988 143664
rect 13748 2128 14988 143664
rect 23748 2128 24988 143664
rect 33748 2128 34988 143664
rect 43748 2128 44988 143664
rect 53748 2128 54988 143664
rect 63748 2128 64988 143664
rect 73748 2128 74988 143664
rect 83748 2128 84988 143664
rect 93748 2128 94988 143664
rect 103748 2128 104988 143664
rect 113748 2128 114988 143664
rect 123748 2128 124988 143664
rect 133748 2128 134988 143664
<< obsm4 >>
rect 9627 2483 13668 143445
rect 15068 2483 23668 143445
rect 25068 2483 33668 143445
rect 35068 2483 43668 143445
rect 45068 2483 53668 143445
rect 55068 2483 63668 143445
rect 65068 2483 73668 143445
rect 75068 2483 83668 143445
rect 85068 2483 93668 143445
rect 95068 2483 103668 143445
rect 105068 2483 113668 143445
rect 115068 2483 123668 143445
rect 125068 2483 133668 143445
rect 135068 2483 141989 143445
<< labels >>
rlabel metal3 s 142965 5720 143765 5840 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 140042 145109 140098 145909 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 124310 145109 124366 145909 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 108578 145109 108634 145909 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 92846 145109 92902 145909 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 77114 145109 77170 145909 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 61382 145109 61438 145909 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 45650 145109 45706 145909 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 29918 145109 29974 145909 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 14186 145109 14242 145909 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 142965 19592 143765 19712 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 134104 800 134224 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 126760 800 126880 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 112072 800 112192 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 142965 33464 143765 33584 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 142965 47336 143765 47456 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 142965 61208 143765 61328 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 142965 75080 143765 75200 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 142965 88952 143765 89072 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 142965 102824 143765 102944 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 142965 116696 143765 116816 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 142965 130568 143765 130688 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 142965 14968 143765 15088 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 129554 145109 129610 145909 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 113822 145109 113878 145909 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 98090 145109 98146 145909 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 82358 145109 82414 145909 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 66626 145109 66682 145909 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 50894 145109 50950 145909 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 35162 145109 35218 145909 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 19430 145109 19486 145909 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 3698 145109 3754 145909 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 136552 800 136672 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 142965 28840 143765 28960 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 0 121864 800 121984 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 114520 800 114640 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 0 107176 800 107296 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 77800 800 77920 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 142965 42712 143765 42832 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 142965 56584 143765 56704 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 142965 70456 143765 70576 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 142965 84328 143765 84448 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 142965 98200 143765 98320 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 142965 112072 143765 112192 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 142965 125944 143765 126064 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 142965 139816 143765 139936 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 142965 10344 143765 10464 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 134798 145109 134854 145909 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 119066 145109 119122 145909 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 103334 145109 103390 145909 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 87602 145109 87658 145909 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 71870 145109 71926 145909 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 56138 145109 56194 145909 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 40406 145109 40462 145909 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 24674 145109 24730 145909 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 8942 145109 8998 145909 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 142965 24216 143765 24336 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 0 131656 800 131776 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 124312 800 124432 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 0 109624 800 109744 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 142965 38088 143765 38208 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 142965 51960 143765 52080 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 142965 65832 143765 65952 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 142965 79704 143765 79824 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 142965 93576 143765 93696 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 142965 107448 143765 107568 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 142965 121320 143765 121440 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 142965 135192 143765 135312 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 139214 0 139270 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 134522 0 134578 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 135350 0 135406 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 136178 0 136234 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 137006 0 137062 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 138662 0 138718 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 99746 0 99802 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 107198 0 107254 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 3748 2128 4988 143664 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 23748 2128 24988 143664 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 43748 2128 44988 143664 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 63748 2128 64988 143664 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 83748 2128 84988 143664 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 103748 2128 104988 143664 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 123748 2128 124988 143664 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 13748 2128 14988 143664 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 33748 2128 34988 143664 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 53748 2128 54988 143664 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 73748 2128 74988 143664 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 93748 2128 94988 143664 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 113748 2128 114988 143664 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 133748 2128 134988 143664 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 3974 0 4030 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 143765 145909
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 70062540
string GDS_FILE /home/ejjimenezu/Repos/caravel_simple_fpu/openlane/fpu/runs/24_12_04_06_36/results/signoff/fpu.magic.gds
string GDS_START 1102790
<< end >>

