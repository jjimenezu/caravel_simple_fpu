magic
tech sky130A
magscale 1 2
timestamp 1733361216
<< obsli1 >>
rect 1104 2159 174248 175185
<< obsm1 >>
rect 934 1232 174248 175216
<< metal2 >>
rect 3882 176698 3938 177498
rect 10322 176698 10378 177498
rect 16762 176698 16818 177498
rect 23202 176698 23258 177498
rect 29642 176698 29698 177498
rect 36082 176698 36138 177498
rect 42522 176698 42578 177498
rect 48962 176698 49018 177498
rect 55402 176698 55458 177498
rect 61842 176698 61898 177498
rect 68282 176698 68338 177498
rect 74722 176698 74778 177498
rect 81162 176698 81218 177498
rect 87602 176698 87658 177498
rect 94042 176698 94098 177498
rect 100482 176698 100538 177498
rect 106922 176698 106978 177498
rect 113362 176698 113418 177498
rect 119802 176698 119858 177498
rect 126242 176698 126298 177498
rect 132682 176698 132738 177498
rect 139122 176698 139178 177498
rect 145562 176698 145618 177498
rect 152002 176698 152058 177498
rect 158442 176698 158498 177498
rect 164882 176698 164938 177498
rect 171322 176698 171378 177498
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54758 0 54814 800
rect 55034 0 55090 800
rect 55310 0 55366 800
rect 55586 0 55642 800
rect 55862 0 55918 800
rect 56138 0 56194 800
rect 56414 0 56470 800
rect 56690 0 56746 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58622 0 58678 800
rect 58898 0 58954 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59726 0 59782 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61382 0 61438 800
rect 61658 0 61714 800
rect 61934 0 61990 800
rect 62210 0 62266 800
rect 62486 0 62542 800
rect 62762 0 62818 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63590 0 63646 800
rect 63866 0 63922 800
rect 64142 0 64198 800
rect 64418 0 64474 800
rect 64694 0 64750 800
rect 64970 0 65026 800
rect 65246 0 65302 800
rect 65522 0 65578 800
rect 65798 0 65854 800
rect 66074 0 66130 800
rect 66350 0 66406 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 68006 0 68062 800
rect 68282 0 68338 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69110 0 69166 800
rect 69386 0 69442 800
rect 69662 0 69718 800
rect 69938 0 69994 800
rect 70214 0 70270 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 71042 0 71098 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71870 0 71926 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72698 0 72754 800
rect 72974 0 73030 800
rect 73250 0 73306 800
rect 73526 0 73582 800
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75182 0 75238 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 76010 0 76066 800
rect 76286 0 76342 800
rect 76562 0 76618 800
rect 76838 0 76894 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78770 0 78826 800
rect 79046 0 79102 800
rect 79322 0 79378 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80150 0 80206 800
rect 80426 0 80482 800
rect 80702 0 80758 800
rect 80978 0 81034 800
rect 81254 0 81310 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 82082 0 82138 800
rect 82358 0 82414 800
rect 82634 0 82690 800
rect 82910 0 82966 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83738 0 83794 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84566 0 84622 800
rect 84842 0 84898 800
rect 85118 0 85174 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 85946 0 86002 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86774 0 86830 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87602 0 87658 800
rect 87878 0 87934 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88706 0 88762 800
rect 88982 0 89038 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89810 0 89866 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90638 0 90694 800
rect 90914 0 90970 800
rect 91190 0 91246 800
rect 91466 0 91522 800
rect 91742 0 91798 800
rect 92018 0 92074 800
rect 92294 0 92350 800
rect 92570 0 92626 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93674 0 93730 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94502 0 94558 800
rect 94778 0 94834 800
rect 95054 0 95110 800
rect 95330 0 95386 800
rect 95606 0 95662 800
rect 95882 0 95938 800
rect 96158 0 96214 800
rect 96434 0 96490 800
rect 96710 0 96766 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97538 0 97594 800
rect 97814 0 97870 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99194 0 99250 800
rect 99470 0 99526 800
rect 99746 0 99802 800
rect 100022 0 100078 800
rect 100298 0 100354 800
rect 100574 0 100630 800
rect 100850 0 100906 800
rect 101126 0 101182 800
rect 101402 0 101458 800
rect 101678 0 101734 800
rect 101954 0 102010 800
rect 102230 0 102286 800
rect 102506 0 102562 800
rect 102782 0 102838 800
rect 103058 0 103114 800
rect 103334 0 103390 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104714 0 104770 800
rect 104990 0 105046 800
rect 105266 0 105322 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106094 0 106150 800
rect 106370 0 106426 800
rect 106646 0 106702 800
rect 106922 0 106978 800
rect 107198 0 107254 800
rect 107474 0 107530 800
rect 107750 0 107806 800
rect 108026 0 108082 800
rect 108302 0 108358 800
rect 108578 0 108634 800
rect 108854 0 108910 800
rect 109130 0 109186 800
rect 109406 0 109462 800
rect 109682 0 109738 800
rect 109958 0 110014 800
rect 110234 0 110290 800
rect 110510 0 110566 800
rect 110786 0 110842 800
rect 111062 0 111118 800
rect 111338 0 111394 800
rect 111614 0 111670 800
rect 111890 0 111946 800
rect 112166 0 112222 800
rect 112442 0 112498 800
rect 112718 0 112774 800
rect 112994 0 113050 800
rect 113270 0 113326 800
rect 113546 0 113602 800
rect 113822 0 113878 800
rect 114098 0 114154 800
rect 114374 0 114430 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115202 0 115258 800
rect 115478 0 115534 800
rect 115754 0 115810 800
rect 116030 0 116086 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117134 0 117190 800
rect 117410 0 117466 800
rect 117686 0 117742 800
rect 117962 0 118018 800
rect 118238 0 118294 800
rect 118514 0 118570 800
rect 118790 0 118846 800
rect 119066 0 119122 800
rect 119342 0 119398 800
rect 119618 0 119674 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120446 0 120502 800
rect 120722 0 120778 800
rect 120998 0 121054 800
rect 121274 0 121330 800
rect 121550 0 121606 800
rect 121826 0 121882 800
rect 122102 0 122158 800
rect 122378 0 122434 800
rect 122654 0 122710 800
rect 122930 0 122986 800
rect 123206 0 123262 800
rect 123482 0 123538 800
rect 123758 0 123814 800
rect 124034 0 124090 800
rect 124310 0 124366 800
rect 124586 0 124642 800
rect 124862 0 124918 800
rect 125138 0 125194 800
rect 125414 0 125470 800
rect 125690 0 125746 800
rect 125966 0 126022 800
rect 126242 0 126298 800
rect 126518 0 126574 800
rect 126794 0 126850 800
rect 127070 0 127126 800
rect 127346 0 127402 800
rect 127622 0 127678 800
rect 127898 0 127954 800
rect 128174 0 128230 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129002 0 129058 800
rect 129278 0 129334 800
rect 129554 0 129610 800
rect 129830 0 129886 800
rect 130106 0 130162 800
rect 130382 0 130438 800
rect 130658 0 130714 800
rect 130934 0 130990 800
rect 131210 0 131266 800
rect 131486 0 131542 800
rect 131762 0 131818 800
rect 132038 0 132094 800
rect 132314 0 132370 800
rect 132590 0 132646 800
rect 132866 0 132922 800
rect 133142 0 133198 800
rect 133418 0 133474 800
rect 133694 0 133750 800
rect 133970 0 134026 800
rect 134246 0 134302 800
rect 134522 0 134578 800
rect 134798 0 134854 800
rect 135074 0 135130 800
rect 135350 0 135406 800
rect 135626 0 135682 800
rect 135902 0 135958 800
rect 136178 0 136234 800
rect 136454 0 136510 800
rect 136730 0 136786 800
rect 137006 0 137062 800
rect 137282 0 137338 800
rect 137558 0 137614 800
rect 137834 0 137890 800
rect 138110 0 138166 800
rect 138386 0 138442 800
rect 138662 0 138718 800
rect 138938 0 138994 800
rect 139214 0 139270 800
rect 139490 0 139546 800
rect 139766 0 139822 800
rect 140042 0 140098 800
rect 140318 0 140374 800
rect 140594 0 140650 800
rect 140870 0 140926 800
rect 141146 0 141202 800
rect 141422 0 141478 800
rect 141698 0 141754 800
rect 141974 0 142030 800
rect 142250 0 142306 800
rect 142526 0 142582 800
rect 142802 0 142858 800
rect 143078 0 143134 800
rect 143354 0 143410 800
rect 143630 0 143686 800
rect 143906 0 143962 800
rect 144182 0 144238 800
rect 144458 0 144514 800
rect 144734 0 144790 800
rect 145010 0 145066 800
rect 145286 0 145342 800
rect 145562 0 145618 800
rect 145838 0 145894 800
rect 146114 0 146170 800
rect 146390 0 146446 800
rect 146666 0 146722 800
rect 146942 0 146998 800
rect 147218 0 147274 800
rect 147494 0 147550 800
rect 147770 0 147826 800
rect 148046 0 148102 800
rect 148322 0 148378 800
rect 148598 0 148654 800
rect 148874 0 148930 800
rect 149150 0 149206 800
rect 149426 0 149482 800
rect 149702 0 149758 800
rect 149978 0 150034 800
rect 150254 0 150310 800
rect 150530 0 150586 800
rect 150806 0 150862 800
rect 151082 0 151138 800
rect 151358 0 151414 800
rect 151634 0 151690 800
rect 151910 0 151966 800
rect 152186 0 152242 800
rect 152462 0 152518 800
rect 152738 0 152794 800
rect 153014 0 153070 800
rect 153290 0 153346 800
rect 153566 0 153622 800
rect 153842 0 153898 800
rect 154118 0 154174 800
rect 154394 0 154450 800
rect 154670 0 154726 800
rect 154946 0 155002 800
rect 155222 0 155278 800
rect 155498 0 155554 800
<< obsm2 >>
rect 938 176642 3826 176746
rect 3994 176642 10266 176746
rect 10434 176642 16706 176746
rect 16874 176642 23146 176746
rect 23314 176642 29586 176746
rect 29754 176642 36026 176746
rect 36194 176642 42466 176746
rect 42634 176642 48906 176746
rect 49074 176642 55346 176746
rect 55514 176642 61786 176746
rect 61954 176642 68226 176746
rect 68394 176642 74666 176746
rect 74834 176642 81106 176746
rect 81274 176642 87546 176746
rect 87714 176642 93986 176746
rect 94154 176642 100426 176746
rect 100594 176642 106866 176746
rect 107034 176642 113306 176746
rect 113474 176642 119746 176746
rect 119914 176642 126186 176746
rect 126354 176642 132626 176746
rect 132794 176642 139066 176746
rect 139234 176642 145506 176746
rect 145674 176642 151946 176746
rect 152114 176642 158386 176746
rect 158554 176642 164826 176746
rect 164994 176642 171266 176746
rect 171434 176642 174138 176746
rect 938 856 174138 176642
rect 938 800 19650 856
rect 19818 800 19926 856
rect 20094 800 20202 856
rect 20370 800 20478 856
rect 20646 800 20754 856
rect 20922 800 21030 856
rect 21198 800 21306 856
rect 21474 800 21582 856
rect 21750 800 21858 856
rect 22026 800 22134 856
rect 22302 800 22410 856
rect 22578 800 22686 856
rect 22854 800 22962 856
rect 23130 800 23238 856
rect 23406 800 23514 856
rect 23682 800 23790 856
rect 23958 800 24066 856
rect 24234 800 24342 856
rect 24510 800 24618 856
rect 24786 800 24894 856
rect 25062 800 25170 856
rect 25338 800 25446 856
rect 25614 800 25722 856
rect 25890 800 25998 856
rect 26166 800 26274 856
rect 26442 800 26550 856
rect 26718 800 26826 856
rect 26994 800 27102 856
rect 27270 800 27378 856
rect 27546 800 27654 856
rect 27822 800 27930 856
rect 28098 800 28206 856
rect 28374 800 28482 856
rect 28650 800 28758 856
rect 28926 800 29034 856
rect 29202 800 29310 856
rect 29478 800 29586 856
rect 29754 800 29862 856
rect 30030 800 30138 856
rect 30306 800 30414 856
rect 30582 800 30690 856
rect 30858 800 30966 856
rect 31134 800 31242 856
rect 31410 800 31518 856
rect 31686 800 31794 856
rect 31962 800 32070 856
rect 32238 800 32346 856
rect 32514 800 32622 856
rect 32790 800 32898 856
rect 33066 800 33174 856
rect 33342 800 33450 856
rect 33618 800 33726 856
rect 33894 800 34002 856
rect 34170 800 34278 856
rect 34446 800 34554 856
rect 34722 800 34830 856
rect 34998 800 35106 856
rect 35274 800 35382 856
rect 35550 800 35658 856
rect 35826 800 35934 856
rect 36102 800 36210 856
rect 36378 800 36486 856
rect 36654 800 36762 856
rect 36930 800 37038 856
rect 37206 800 37314 856
rect 37482 800 37590 856
rect 37758 800 37866 856
rect 38034 800 38142 856
rect 38310 800 38418 856
rect 38586 800 38694 856
rect 38862 800 38970 856
rect 39138 800 39246 856
rect 39414 800 39522 856
rect 39690 800 39798 856
rect 39966 800 40074 856
rect 40242 800 40350 856
rect 40518 800 40626 856
rect 40794 800 40902 856
rect 41070 800 41178 856
rect 41346 800 41454 856
rect 41622 800 41730 856
rect 41898 800 42006 856
rect 42174 800 42282 856
rect 42450 800 42558 856
rect 42726 800 42834 856
rect 43002 800 43110 856
rect 43278 800 43386 856
rect 43554 800 43662 856
rect 43830 800 43938 856
rect 44106 800 44214 856
rect 44382 800 44490 856
rect 44658 800 44766 856
rect 44934 800 45042 856
rect 45210 800 45318 856
rect 45486 800 45594 856
rect 45762 800 45870 856
rect 46038 800 46146 856
rect 46314 800 46422 856
rect 46590 800 46698 856
rect 46866 800 46974 856
rect 47142 800 47250 856
rect 47418 800 47526 856
rect 47694 800 47802 856
rect 47970 800 48078 856
rect 48246 800 48354 856
rect 48522 800 48630 856
rect 48798 800 48906 856
rect 49074 800 49182 856
rect 49350 800 49458 856
rect 49626 800 49734 856
rect 49902 800 50010 856
rect 50178 800 50286 856
rect 50454 800 50562 856
rect 50730 800 50838 856
rect 51006 800 51114 856
rect 51282 800 51390 856
rect 51558 800 51666 856
rect 51834 800 51942 856
rect 52110 800 52218 856
rect 52386 800 52494 856
rect 52662 800 52770 856
rect 52938 800 53046 856
rect 53214 800 53322 856
rect 53490 800 53598 856
rect 53766 800 53874 856
rect 54042 800 54150 856
rect 54318 800 54426 856
rect 54594 800 54702 856
rect 54870 800 54978 856
rect 55146 800 55254 856
rect 55422 800 55530 856
rect 55698 800 55806 856
rect 55974 800 56082 856
rect 56250 800 56358 856
rect 56526 800 56634 856
rect 56802 800 56910 856
rect 57078 800 57186 856
rect 57354 800 57462 856
rect 57630 800 57738 856
rect 57906 800 58014 856
rect 58182 800 58290 856
rect 58458 800 58566 856
rect 58734 800 58842 856
rect 59010 800 59118 856
rect 59286 800 59394 856
rect 59562 800 59670 856
rect 59838 800 59946 856
rect 60114 800 60222 856
rect 60390 800 60498 856
rect 60666 800 60774 856
rect 60942 800 61050 856
rect 61218 800 61326 856
rect 61494 800 61602 856
rect 61770 800 61878 856
rect 62046 800 62154 856
rect 62322 800 62430 856
rect 62598 800 62706 856
rect 62874 800 62982 856
rect 63150 800 63258 856
rect 63426 800 63534 856
rect 63702 800 63810 856
rect 63978 800 64086 856
rect 64254 800 64362 856
rect 64530 800 64638 856
rect 64806 800 64914 856
rect 65082 800 65190 856
rect 65358 800 65466 856
rect 65634 800 65742 856
rect 65910 800 66018 856
rect 66186 800 66294 856
rect 66462 800 66570 856
rect 66738 800 66846 856
rect 67014 800 67122 856
rect 67290 800 67398 856
rect 67566 800 67674 856
rect 67842 800 67950 856
rect 68118 800 68226 856
rect 68394 800 68502 856
rect 68670 800 68778 856
rect 68946 800 69054 856
rect 69222 800 69330 856
rect 69498 800 69606 856
rect 69774 800 69882 856
rect 70050 800 70158 856
rect 70326 800 70434 856
rect 70602 800 70710 856
rect 70878 800 70986 856
rect 71154 800 71262 856
rect 71430 800 71538 856
rect 71706 800 71814 856
rect 71982 800 72090 856
rect 72258 800 72366 856
rect 72534 800 72642 856
rect 72810 800 72918 856
rect 73086 800 73194 856
rect 73362 800 73470 856
rect 73638 800 73746 856
rect 73914 800 74022 856
rect 74190 800 74298 856
rect 74466 800 74574 856
rect 74742 800 74850 856
rect 75018 800 75126 856
rect 75294 800 75402 856
rect 75570 800 75678 856
rect 75846 800 75954 856
rect 76122 800 76230 856
rect 76398 800 76506 856
rect 76674 800 76782 856
rect 76950 800 77058 856
rect 77226 800 77334 856
rect 77502 800 77610 856
rect 77778 800 77886 856
rect 78054 800 78162 856
rect 78330 800 78438 856
rect 78606 800 78714 856
rect 78882 800 78990 856
rect 79158 800 79266 856
rect 79434 800 79542 856
rect 79710 800 79818 856
rect 79986 800 80094 856
rect 80262 800 80370 856
rect 80538 800 80646 856
rect 80814 800 80922 856
rect 81090 800 81198 856
rect 81366 800 81474 856
rect 81642 800 81750 856
rect 81918 800 82026 856
rect 82194 800 82302 856
rect 82470 800 82578 856
rect 82746 800 82854 856
rect 83022 800 83130 856
rect 83298 800 83406 856
rect 83574 800 83682 856
rect 83850 800 83958 856
rect 84126 800 84234 856
rect 84402 800 84510 856
rect 84678 800 84786 856
rect 84954 800 85062 856
rect 85230 800 85338 856
rect 85506 800 85614 856
rect 85782 800 85890 856
rect 86058 800 86166 856
rect 86334 800 86442 856
rect 86610 800 86718 856
rect 86886 800 86994 856
rect 87162 800 87270 856
rect 87438 800 87546 856
rect 87714 800 87822 856
rect 87990 800 88098 856
rect 88266 800 88374 856
rect 88542 800 88650 856
rect 88818 800 88926 856
rect 89094 800 89202 856
rect 89370 800 89478 856
rect 89646 800 89754 856
rect 89922 800 90030 856
rect 90198 800 90306 856
rect 90474 800 90582 856
rect 90750 800 90858 856
rect 91026 800 91134 856
rect 91302 800 91410 856
rect 91578 800 91686 856
rect 91854 800 91962 856
rect 92130 800 92238 856
rect 92406 800 92514 856
rect 92682 800 92790 856
rect 92958 800 93066 856
rect 93234 800 93342 856
rect 93510 800 93618 856
rect 93786 800 93894 856
rect 94062 800 94170 856
rect 94338 800 94446 856
rect 94614 800 94722 856
rect 94890 800 94998 856
rect 95166 800 95274 856
rect 95442 800 95550 856
rect 95718 800 95826 856
rect 95994 800 96102 856
rect 96270 800 96378 856
rect 96546 800 96654 856
rect 96822 800 96930 856
rect 97098 800 97206 856
rect 97374 800 97482 856
rect 97650 800 97758 856
rect 97926 800 98034 856
rect 98202 800 98310 856
rect 98478 800 98586 856
rect 98754 800 98862 856
rect 99030 800 99138 856
rect 99306 800 99414 856
rect 99582 800 99690 856
rect 99858 800 99966 856
rect 100134 800 100242 856
rect 100410 800 100518 856
rect 100686 800 100794 856
rect 100962 800 101070 856
rect 101238 800 101346 856
rect 101514 800 101622 856
rect 101790 800 101898 856
rect 102066 800 102174 856
rect 102342 800 102450 856
rect 102618 800 102726 856
rect 102894 800 103002 856
rect 103170 800 103278 856
rect 103446 800 103554 856
rect 103722 800 103830 856
rect 103998 800 104106 856
rect 104274 800 104382 856
rect 104550 800 104658 856
rect 104826 800 104934 856
rect 105102 800 105210 856
rect 105378 800 105486 856
rect 105654 800 105762 856
rect 105930 800 106038 856
rect 106206 800 106314 856
rect 106482 800 106590 856
rect 106758 800 106866 856
rect 107034 800 107142 856
rect 107310 800 107418 856
rect 107586 800 107694 856
rect 107862 800 107970 856
rect 108138 800 108246 856
rect 108414 800 108522 856
rect 108690 800 108798 856
rect 108966 800 109074 856
rect 109242 800 109350 856
rect 109518 800 109626 856
rect 109794 800 109902 856
rect 110070 800 110178 856
rect 110346 800 110454 856
rect 110622 800 110730 856
rect 110898 800 111006 856
rect 111174 800 111282 856
rect 111450 800 111558 856
rect 111726 800 111834 856
rect 112002 800 112110 856
rect 112278 800 112386 856
rect 112554 800 112662 856
rect 112830 800 112938 856
rect 113106 800 113214 856
rect 113382 800 113490 856
rect 113658 800 113766 856
rect 113934 800 114042 856
rect 114210 800 114318 856
rect 114486 800 114594 856
rect 114762 800 114870 856
rect 115038 800 115146 856
rect 115314 800 115422 856
rect 115590 800 115698 856
rect 115866 800 115974 856
rect 116142 800 116250 856
rect 116418 800 116526 856
rect 116694 800 116802 856
rect 116970 800 117078 856
rect 117246 800 117354 856
rect 117522 800 117630 856
rect 117798 800 117906 856
rect 118074 800 118182 856
rect 118350 800 118458 856
rect 118626 800 118734 856
rect 118902 800 119010 856
rect 119178 800 119286 856
rect 119454 800 119562 856
rect 119730 800 119838 856
rect 120006 800 120114 856
rect 120282 800 120390 856
rect 120558 800 120666 856
rect 120834 800 120942 856
rect 121110 800 121218 856
rect 121386 800 121494 856
rect 121662 800 121770 856
rect 121938 800 122046 856
rect 122214 800 122322 856
rect 122490 800 122598 856
rect 122766 800 122874 856
rect 123042 800 123150 856
rect 123318 800 123426 856
rect 123594 800 123702 856
rect 123870 800 123978 856
rect 124146 800 124254 856
rect 124422 800 124530 856
rect 124698 800 124806 856
rect 124974 800 125082 856
rect 125250 800 125358 856
rect 125526 800 125634 856
rect 125802 800 125910 856
rect 126078 800 126186 856
rect 126354 800 126462 856
rect 126630 800 126738 856
rect 126906 800 127014 856
rect 127182 800 127290 856
rect 127458 800 127566 856
rect 127734 800 127842 856
rect 128010 800 128118 856
rect 128286 800 128394 856
rect 128562 800 128670 856
rect 128838 800 128946 856
rect 129114 800 129222 856
rect 129390 800 129498 856
rect 129666 800 129774 856
rect 129942 800 130050 856
rect 130218 800 130326 856
rect 130494 800 130602 856
rect 130770 800 130878 856
rect 131046 800 131154 856
rect 131322 800 131430 856
rect 131598 800 131706 856
rect 131874 800 131982 856
rect 132150 800 132258 856
rect 132426 800 132534 856
rect 132702 800 132810 856
rect 132978 800 133086 856
rect 133254 800 133362 856
rect 133530 800 133638 856
rect 133806 800 133914 856
rect 134082 800 134190 856
rect 134358 800 134466 856
rect 134634 800 134742 856
rect 134910 800 135018 856
rect 135186 800 135294 856
rect 135462 800 135570 856
rect 135738 800 135846 856
rect 136014 800 136122 856
rect 136290 800 136398 856
rect 136566 800 136674 856
rect 136842 800 136950 856
rect 137118 800 137226 856
rect 137394 800 137502 856
rect 137670 800 137778 856
rect 137946 800 138054 856
rect 138222 800 138330 856
rect 138498 800 138606 856
rect 138774 800 138882 856
rect 139050 800 139158 856
rect 139326 800 139434 856
rect 139602 800 139710 856
rect 139878 800 139986 856
rect 140154 800 140262 856
rect 140430 800 140538 856
rect 140706 800 140814 856
rect 140982 800 141090 856
rect 141258 800 141366 856
rect 141534 800 141642 856
rect 141810 800 141918 856
rect 142086 800 142194 856
rect 142362 800 142470 856
rect 142638 800 142746 856
rect 142914 800 143022 856
rect 143190 800 143298 856
rect 143466 800 143574 856
rect 143742 800 143850 856
rect 144018 800 144126 856
rect 144294 800 144402 856
rect 144570 800 144678 856
rect 144846 800 144954 856
rect 145122 800 145230 856
rect 145398 800 145506 856
rect 145674 800 145782 856
rect 145950 800 146058 856
rect 146226 800 146334 856
rect 146502 800 146610 856
rect 146778 800 146886 856
rect 147054 800 147162 856
rect 147330 800 147438 856
rect 147606 800 147714 856
rect 147882 800 147990 856
rect 148158 800 148266 856
rect 148434 800 148542 856
rect 148710 800 148818 856
rect 148986 800 149094 856
rect 149262 800 149370 856
rect 149538 800 149646 856
rect 149814 800 149922 856
rect 150090 800 150198 856
rect 150366 800 150474 856
rect 150642 800 150750 856
rect 150918 800 151026 856
rect 151194 800 151302 856
rect 151470 800 151578 856
rect 151746 800 151854 856
rect 152022 800 152130 856
rect 152298 800 152406 856
rect 152574 800 152682 856
rect 152850 800 152958 856
rect 153126 800 153234 856
rect 153402 800 153510 856
rect 153678 800 153786 856
rect 153954 800 154062 856
rect 154230 800 154338 856
rect 154506 800 154614 856
rect 154782 800 154890 856
rect 155058 800 155166 856
rect 155334 800 155442 856
rect 155610 800 174138 856
<< metal3 >>
rect 0 172456 800 172576
rect 174554 171368 175354 171488
rect 0 169464 800 169584
rect 0 166472 800 166592
rect 174554 165656 175354 165776
rect 0 163480 800 163600
rect 0 160488 800 160608
rect 174554 159944 175354 160064
rect 0 157496 800 157616
rect 0 154504 800 154624
rect 174554 154232 175354 154352
rect 0 151512 800 151632
rect 0 148520 800 148640
rect 174554 148520 175354 148640
rect 0 145528 800 145648
rect 174554 142808 175354 142928
rect 0 142536 800 142656
rect 0 139544 800 139664
rect 174554 137096 175354 137216
rect 0 136552 800 136672
rect 0 133560 800 133680
rect 174554 131384 175354 131504
rect 0 130568 800 130688
rect 0 127576 800 127696
rect 174554 125672 175354 125792
rect 0 124584 800 124704
rect 0 121592 800 121712
rect 174554 119960 175354 120080
rect 0 118600 800 118720
rect 0 115608 800 115728
rect 174554 114248 175354 114368
rect 0 112616 800 112736
rect 0 109624 800 109744
rect 174554 108536 175354 108656
rect 0 106632 800 106752
rect 0 103640 800 103760
rect 174554 102824 175354 102944
rect 0 100648 800 100768
rect 0 97656 800 97776
rect 174554 97112 175354 97232
rect 0 94664 800 94784
rect 0 91672 800 91792
rect 174554 91400 175354 91520
rect 0 88680 800 88800
rect 0 85688 800 85808
rect 174554 85688 175354 85808
rect 0 82696 800 82816
rect 174554 79976 175354 80096
rect 0 79704 800 79824
rect 0 76712 800 76832
rect 174554 74264 175354 74384
rect 0 73720 800 73840
rect 0 70728 800 70848
rect 174554 68552 175354 68672
rect 0 67736 800 67856
rect 0 64744 800 64864
rect 174554 62840 175354 62960
rect 0 61752 800 61872
rect 0 58760 800 58880
rect 174554 57128 175354 57248
rect 0 55768 800 55888
rect 0 52776 800 52896
rect 174554 51416 175354 51536
rect 0 49784 800 49904
rect 0 46792 800 46912
rect 174554 45704 175354 45824
rect 0 43800 800 43920
rect 0 40808 800 40928
rect 174554 39992 175354 40112
rect 0 37816 800 37936
rect 0 34824 800 34944
rect 174554 34280 175354 34400
rect 0 31832 800 31952
rect 0 28840 800 28960
rect 174554 28568 175354 28688
rect 0 25848 800 25968
rect 0 22856 800 22976
rect 174554 22856 175354 22976
rect 0 19864 800 19984
rect 174554 17144 175354 17264
rect 0 16872 800 16992
rect 0 13880 800 14000
rect 174554 11432 175354 11552
rect 0 10888 800 11008
rect 0 7896 800 8016
rect 174554 5720 175354 5840
rect 0 4904 800 5024
<< obsm3 >>
rect 798 172656 174554 175201
rect 880 172376 174554 172656
rect 798 171568 174554 172376
rect 798 171288 174474 171568
rect 798 169664 174554 171288
rect 880 169384 174554 169664
rect 798 166672 174554 169384
rect 880 166392 174554 166672
rect 798 165856 174554 166392
rect 798 165576 174474 165856
rect 798 163680 174554 165576
rect 880 163400 174554 163680
rect 798 160688 174554 163400
rect 880 160408 174554 160688
rect 798 160144 174554 160408
rect 798 159864 174474 160144
rect 798 157696 174554 159864
rect 880 157416 174554 157696
rect 798 154704 174554 157416
rect 880 154432 174554 154704
rect 880 154424 174474 154432
rect 798 154152 174474 154424
rect 798 151712 174554 154152
rect 880 151432 174554 151712
rect 798 148720 174554 151432
rect 880 148440 174474 148720
rect 798 145728 174554 148440
rect 880 145448 174554 145728
rect 798 143008 174554 145448
rect 798 142736 174474 143008
rect 880 142728 174474 142736
rect 880 142456 174554 142728
rect 798 139744 174554 142456
rect 880 139464 174554 139744
rect 798 137296 174554 139464
rect 798 137016 174474 137296
rect 798 136752 174554 137016
rect 880 136472 174554 136752
rect 798 133760 174554 136472
rect 880 133480 174554 133760
rect 798 131584 174554 133480
rect 798 131304 174474 131584
rect 798 130768 174554 131304
rect 880 130488 174554 130768
rect 798 127776 174554 130488
rect 880 127496 174554 127776
rect 798 125872 174554 127496
rect 798 125592 174474 125872
rect 798 124784 174554 125592
rect 880 124504 174554 124784
rect 798 121792 174554 124504
rect 880 121512 174554 121792
rect 798 120160 174554 121512
rect 798 119880 174474 120160
rect 798 118800 174554 119880
rect 880 118520 174554 118800
rect 798 115808 174554 118520
rect 880 115528 174554 115808
rect 798 114448 174554 115528
rect 798 114168 174474 114448
rect 798 112816 174554 114168
rect 880 112536 174554 112816
rect 798 109824 174554 112536
rect 880 109544 174554 109824
rect 798 108736 174554 109544
rect 798 108456 174474 108736
rect 798 106832 174554 108456
rect 880 106552 174554 106832
rect 798 103840 174554 106552
rect 880 103560 174554 103840
rect 798 103024 174554 103560
rect 798 102744 174474 103024
rect 798 100848 174554 102744
rect 880 100568 174554 100848
rect 798 97856 174554 100568
rect 880 97576 174554 97856
rect 798 97312 174554 97576
rect 798 97032 174474 97312
rect 798 94864 174554 97032
rect 880 94584 174554 94864
rect 798 91872 174554 94584
rect 880 91600 174554 91872
rect 880 91592 174474 91600
rect 798 91320 174474 91592
rect 798 88880 174554 91320
rect 880 88600 174554 88880
rect 798 85888 174554 88600
rect 880 85608 174474 85888
rect 798 82896 174554 85608
rect 880 82616 174554 82896
rect 798 80176 174554 82616
rect 798 79904 174474 80176
rect 880 79896 174474 79904
rect 880 79624 174554 79896
rect 798 76912 174554 79624
rect 880 76632 174554 76912
rect 798 74464 174554 76632
rect 798 74184 174474 74464
rect 798 73920 174554 74184
rect 880 73640 174554 73920
rect 798 70928 174554 73640
rect 880 70648 174554 70928
rect 798 68752 174554 70648
rect 798 68472 174474 68752
rect 798 67936 174554 68472
rect 880 67656 174554 67936
rect 798 64944 174554 67656
rect 880 64664 174554 64944
rect 798 63040 174554 64664
rect 798 62760 174474 63040
rect 798 61952 174554 62760
rect 880 61672 174554 61952
rect 798 58960 174554 61672
rect 880 58680 174554 58960
rect 798 57328 174554 58680
rect 798 57048 174474 57328
rect 798 55968 174554 57048
rect 880 55688 174554 55968
rect 798 52976 174554 55688
rect 880 52696 174554 52976
rect 798 51616 174554 52696
rect 798 51336 174474 51616
rect 798 49984 174554 51336
rect 880 49704 174554 49984
rect 798 46992 174554 49704
rect 880 46712 174554 46992
rect 798 45904 174554 46712
rect 798 45624 174474 45904
rect 798 44000 174554 45624
rect 880 43720 174554 44000
rect 798 41008 174554 43720
rect 880 40728 174554 41008
rect 798 40192 174554 40728
rect 798 39912 174474 40192
rect 798 38016 174554 39912
rect 880 37736 174554 38016
rect 798 35024 174554 37736
rect 880 34744 174554 35024
rect 798 34480 174554 34744
rect 798 34200 174474 34480
rect 798 32032 174554 34200
rect 880 31752 174554 32032
rect 798 29040 174554 31752
rect 880 28768 174554 29040
rect 880 28760 174474 28768
rect 798 28488 174474 28760
rect 798 26048 174554 28488
rect 880 25768 174554 26048
rect 798 23056 174554 25768
rect 880 22776 174474 23056
rect 798 20064 174554 22776
rect 880 19784 174554 20064
rect 798 17344 174554 19784
rect 798 17072 174474 17344
rect 880 17064 174474 17072
rect 880 16792 174554 17064
rect 798 14080 174554 16792
rect 880 13800 174554 14080
rect 798 11632 174554 13800
rect 798 11352 174474 11632
rect 798 11088 174554 11352
rect 880 10808 174554 11088
rect 798 8096 174554 10808
rect 880 7816 174554 8096
rect 798 5920 174554 7816
rect 798 5640 174474 5920
rect 798 5104 174554 5640
rect 880 4824 174554 5104
rect 798 1667 174554 4824
<< metal4 >>
rect 3748 2128 4988 175216
rect 13748 2128 14988 175216
rect 23748 2128 24988 175216
rect 33748 2128 34988 175216
rect 43748 2128 44988 175216
rect 53748 2128 54988 175216
rect 63748 2128 64988 175216
rect 73748 2128 74988 175216
rect 83748 2128 84988 175216
rect 93748 2128 94988 175216
rect 103748 2128 104988 175216
rect 113748 2128 114988 175216
rect 123748 2128 124988 175216
rect 133748 2128 134988 175216
rect 143748 2128 144988 175216
rect 153748 2128 154988 175216
rect 163748 2128 164988 175216
<< obsm4 >>
rect 21955 2048 23668 174997
rect 25068 2048 33668 174997
rect 35068 2048 43668 174997
rect 45068 2048 53668 174997
rect 55068 2048 63668 174997
rect 65068 2048 73668 174997
rect 75068 2048 83668 174997
rect 85068 2048 93668 174997
rect 95068 2048 103668 174997
rect 105068 2048 113668 174997
rect 115068 2048 123668 174997
rect 125068 2048 133668 174997
rect 135068 2048 143668 174997
rect 145068 2048 153668 174997
rect 155068 2048 163668 174997
rect 165068 2048 173821 174997
rect 21955 1667 173821 2048
<< labels >>
rlabel metal3 s 174554 5720 175354 5840 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 171322 176698 171378 177498 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 152002 176698 152058 177498 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 132682 176698 132738 177498 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 113362 176698 113418 177498 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 94042 176698 94098 177498 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 74722 176698 74778 177498 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 55402 176698 55458 177498 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 36082 176698 36138 177498 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 16762 176698 16818 177498 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 172456 800 172576 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 174554 22856 175354 22976 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 163480 800 163600 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 154504 800 154624 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 145528 800 145648 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 127576 800 127696 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 118600 800 118720 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 174554 39992 175354 40112 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 174554 57128 175354 57248 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 174554 74264 175354 74384 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 174554 91400 175354 91520 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 174554 108536 175354 108656 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 174554 125672 175354 125792 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 174554 142808 175354 142928 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 174554 159944 175354 160064 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 174554 17144 175354 17264 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 158442 176698 158498 177498 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 139122 176698 139178 177498 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 119802 176698 119858 177498 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 100482 176698 100538 177498 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 81162 176698 81218 177498 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 61842 176698 61898 177498 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 42522 176698 42578 177498 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 23202 176698 23258 177498 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 3882 176698 3938 177498 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 166472 800 166592 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 174554 34280 175354 34400 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 0 157496 800 157616 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 0 148520 800 148640 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 139544 800 139664 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 103640 800 103760 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 94664 800 94784 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 76712 800 76832 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 174554 51416 175354 51536 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 174554 68552 175354 68672 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 174554 85688 175354 85808 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 174554 102824 175354 102944 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 174554 119960 175354 120080 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 174554 137096 175354 137216 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 174554 154232 175354 154352 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 174554 171368 175354 171488 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 174554 11432 175354 11552 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 164882 176698 164938 177498 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 145562 176698 145618 177498 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 126242 176698 126298 177498 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 106922 176698 106978 177498 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 87602 176698 87658 177498 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 68282 176698 68338 177498 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 48962 176698 49018 177498 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 29642 176698 29698 177498 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 10322 176698 10378 177498 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 0 169464 800 169584 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 174554 28568 175354 28688 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 151512 800 151632 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 0 142536 800 142656 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 106632 800 106752 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 88680 800 88800 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 174554 45704 175354 45824 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 174554 62840 175354 62960 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 174554 79976 175354 80096 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 174554 97112 175354 97232 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 174554 114248 175354 114368 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 174554 131384 175354 131504 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 174554 148520 175354 148640 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 174554 165656 175354 165776 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 154946 0 155002 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 134522 0 134578 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 135350 0 135406 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 136178 0 136234 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 137006 0 137062 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 138662 0 138718 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 141146 0 141202 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 142802 0 142858 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 146942 0 146998 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 99746 0 99802 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 107198 0 107254 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 3748 2128 4988 175216 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 23748 2128 24988 175216 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 43748 2128 44988 175216 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 63748 2128 64988 175216 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 83748 2128 84988 175216 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 103748 2128 104988 175216 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 123748 2128 124988 175216 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 143748 2128 144988 175216 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 163748 2128 164988 175216 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 13748 2128 14988 175216 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 33748 2128 34988 175216 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 53748 2128 54988 175216 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 73748 2128 74988 175216 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 93748 2128 94988 175216 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 113748 2128 114988 175216 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 133748 2128 134988 175216 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 153748 2128 154988 175216 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 19706 0 19762 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 175354 177498
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 75407076
string GDS_FILE /home/ejjimenezu/Repos/caravel_simple_fpu/openlane/fpu/runs/24_12_04_18_45/results/signoff/fpu.magic.gds
string GDS_START 1139268
<< end >>

