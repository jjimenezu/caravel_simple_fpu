magic
tech sky130A
magscale 1 2
timestamp 1733402780
<< obsli1 >>
rect 1104 2159 128892 130033
<< obsm1 >>
rect 934 1164 129246 130064
<< metal2 >>
rect 2778 131428 2834 132228
rect 7562 131428 7618 132228
rect 12346 131428 12402 132228
rect 17130 131428 17186 132228
rect 21914 131428 21970 132228
rect 26698 131428 26754 132228
rect 31482 131428 31538 132228
rect 36266 131428 36322 132228
rect 41050 131428 41106 132228
rect 45834 131428 45890 132228
rect 50618 131428 50674 132228
rect 55402 131428 55458 132228
rect 60186 131428 60242 132228
rect 64970 131428 65026 132228
rect 69754 131428 69810 132228
rect 74538 131428 74594 132228
rect 79322 131428 79378 132228
rect 84106 131428 84162 132228
rect 88890 131428 88946 132228
rect 93674 131428 93730 132228
rect 98458 131428 98514 132228
rect 103242 131428 103298 132228
rect 108026 131428 108082 132228
rect 112810 131428 112866 132228
rect 117594 131428 117650 132228
rect 122378 131428 122434 132228
rect 127162 131428 127218 132228
rect 19706 0 19762 800
rect 19890 0 19946 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21730 0 21786 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29642 0 29698 800
rect 29826 0 29882 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31482 0 31538 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34058 0 34114 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36450 0 36506 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 38842 0 38898 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44546 0 44602 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46754 0 46810 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48594 0 48650 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53194 0 53250 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54482 0 54538 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59266 0 59322 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60554 0 60610 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62394 0 62450 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 62946 0 63002 800
rect 63130 0 63186 800
rect 63314 0 63370 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64234 0 64290 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64786 0 64842 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 66074 0 66130 800
rect 66258 0 66314 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68098 0 68154 800
rect 68282 0 68338 800
rect 68466 0 68522 800
rect 68650 0 68706 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 69938 0 69994 800
rect 70122 0 70178 800
rect 70306 0 70362 800
rect 70490 0 70546 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 71962 0 72018 800
rect 72146 0 72202 800
rect 72330 0 72386 800
rect 72514 0 72570 800
rect 72698 0 72754 800
rect 72882 0 72938 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73802 0 73858 800
rect 73986 0 74042 800
rect 74170 0 74226 800
rect 74354 0 74410 800
rect 74538 0 74594 800
rect 74722 0 74778 800
rect 74906 0 74962 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75826 0 75882 800
rect 76010 0 76066 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76562 0 76618 800
rect 76746 0 76802 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77850 0 77906 800
rect 78034 0 78090 800
rect 78218 0 78274 800
rect 78402 0 78458 800
rect 78586 0 78642 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79690 0 79746 800
rect 79874 0 79930 800
rect 80058 0 80114 800
rect 80242 0 80298 800
rect 80426 0 80482 800
rect 80610 0 80666 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82082 0 82138 800
rect 82266 0 82322 800
rect 82450 0 82506 800
rect 82634 0 82690 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83370 0 83426 800
rect 83554 0 83610 800
rect 83738 0 83794 800
rect 83922 0 83978 800
rect 84106 0 84162 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85026 0 85082 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85578 0 85634 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86130 0 86186 800
rect 86314 0 86370 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87418 0 87474 800
rect 87602 0 87658 800
rect 87786 0 87842 800
rect 87970 0 88026 800
rect 88154 0 88210 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89258 0 89314 800
rect 89442 0 89498 800
rect 89626 0 89682 800
rect 89810 0 89866 800
rect 89994 0 90050 800
rect 90178 0 90234 800
rect 90362 0 90418 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91466 0 91522 800
rect 91650 0 91706 800
rect 91834 0 91890 800
rect 92018 0 92074 800
rect 92202 0 92258 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 92938 0 92994 800
rect 93122 0 93178 800
rect 93306 0 93362 800
rect 93490 0 93546 800
rect 93674 0 93730 800
rect 93858 0 93914 800
rect 94042 0 94098 800
rect 94226 0 94282 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95146 0 95202 800
rect 95330 0 95386 800
rect 95514 0 95570 800
rect 95698 0 95754 800
rect 95882 0 95938 800
rect 96066 0 96122 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97170 0 97226 800
rect 97354 0 97410 800
rect 97538 0 97594 800
rect 97722 0 97778 800
rect 97906 0 97962 800
rect 98090 0 98146 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99194 0 99250 800
rect 99378 0 99434 800
rect 99562 0 99618 800
rect 99746 0 99802 800
rect 99930 0 99986 800
rect 100114 0 100170 800
rect 100298 0 100354 800
rect 100482 0 100538 800
rect 100666 0 100722 800
rect 100850 0 100906 800
rect 101034 0 101090 800
rect 101218 0 101274 800
rect 101402 0 101458 800
rect 101586 0 101642 800
rect 101770 0 101826 800
rect 101954 0 102010 800
rect 102138 0 102194 800
rect 102322 0 102378 800
rect 102506 0 102562 800
rect 102690 0 102746 800
rect 102874 0 102930 800
rect 103058 0 103114 800
rect 103242 0 103298 800
rect 103426 0 103482 800
rect 103610 0 103666 800
rect 103794 0 103850 800
rect 103978 0 104034 800
rect 104162 0 104218 800
rect 104346 0 104402 800
rect 104530 0 104586 800
rect 104714 0 104770 800
rect 104898 0 104954 800
rect 105082 0 105138 800
rect 105266 0 105322 800
rect 105450 0 105506 800
rect 105634 0 105690 800
rect 105818 0 105874 800
rect 106002 0 106058 800
rect 106186 0 106242 800
rect 106370 0 106426 800
rect 106554 0 106610 800
rect 106738 0 106794 800
rect 106922 0 106978 800
rect 107106 0 107162 800
rect 107290 0 107346 800
rect 107474 0 107530 800
rect 107658 0 107714 800
rect 107842 0 107898 800
rect 108026 0 108082 800
rect 108210 0 108266 800
rect 108394 0 108450 800
rect 108578 0 108634 800
rect 108762 0 108818 800
rect 108946 0 109002 800
rect 109130 0 109186 800
rect 109314 0 109370 800
rect 109498 0 109554 800
rect 109682 0 109738 800
rect 109866 0 109922 800
rect 110050 0 110106 800
rect 110234 0 110290 800
<< obsm2 >>
rect 938 131372 2722 131458
rect 2890 131372 7506 131458
rect 7674 131372 12290 131458
rect 12458 131372 17074 131458
rect 17242 131372 21858 131458
rect 22026 131372 26642 131458
rect 26810 131372 31426 131458
rect 31594 131372 36210 131458
rect 36378 131372 40994 131458
rect 41162 131372 45778 131458
rect 45946 131372 50562 131458
rect 50730 131372 55346 131458
rect 55514 131372 60130 131458
rect 60298 131372 64914 131458
rect 65082 131372 69698 131458
rect 69866 131372 74482 131458
rect 74650 131372 79266 131458
rect 79434 131372 84050 131458
rect 84218 131372 88834 131458
rect 89002 131372 93618 131458
rect 93786 131372 98402 131458
rect 98570 131372 103186 131458
rect 103354 131372 107970 131458
rect 108138 131372 112754 131458
rect 112922 131372 117538 131458
rect 117706 131372 122322 131458
rect 122490 131372 127106 131458
rect 127274 131372 129240 131458
rect 938 856 129240 131372
rect 938 800 19650 856
rect 19818 800 19834 856
rect 20002 800 20018 856
rect 20186 800 20202 856
rect 20370 800 20386 856
rect 20554 800 20570 856
rect 20738 800 20754 856
rect 20922 800 20938 856
rect 21106 800 21122 856
rect 21290 800 21306 856
rect 21474 800 21490 856
rect 21658 800 21674 856
rect 21842 800 21858 856
rect 22026 800 22042 856
rect 22210 800 22226 856
rect 22394 800 22410 856
rect 22578 800 22594 856
rect 22762 800 22778 856
rect 22946 800 22962 856
rect 23130 800 23146 856
rect 23314 800 23330 856
rect 23498 800 23514 856
rect 23682 800 23698 856
rect 23866 800 23882 856
rect 24050 800 24066 856
rect 24234 800 24250 856
rect 24418 800 24434 856
rect 24602 800 24618 856
rect 24786 800 24802 856
rect 24970 800 24986 856
rect 25154 800 25170 856
rect 25338 800 25354 856
rect 25522 800 25538 856
rect 25706 800 25722 856
rect 25890 800 25906 856
rect 26074 800 26090 856
rect 26258 800 26274 856
rect 26442 800 26458 856
rect 26626 800 26642 856
rect 26810 800 26826 856
rect 26994 800 27010 856
rect 27178 800 27194 856
rect 27362 800 27378 856
rect 27546 800 27562 856
rect 27730 800 27746 856
rect 27914 800 27930 856
rect 28098 800 28114 856
rect 28282 800 28298 856
rect 28466 800 28482 856
rect 28650 800 28666 856
rect 28834 800 28850 856
rect 29018 800 29034 856
rect 29202 800 29218 856
rect 29386 800 29402 856
rect 29570 800 29586 856
rect 29754 800 29770 856
rect 29938 800 29954 856
rect 30122 800 30138 856
rect 30306 800 30322 856
rect 30490 800 30506 856
rect 30674 800 30690 856
rect 30858 800 30874 856
rect 31042 800 31058 856
rect 31226 800 31242 856
rect 31410 800 31426 856
rect 31594 800 31610 856
rect 31778 800 31794 856
rect 31962 800 31978 856
rect 32146 800 32162 856
rect 32330 800 32346 856
rect 32514 800 32530 856
rect 32698 800 32714 856
rect 32882 800 32898 856
rect 33066 800 33082 856
rect 33250 800 33266 856
rect 33434 800 33450 856
rect 33618 800 33634 856
rect 33802 800 33818 856
rect 33986 800 34002 856
rect 34170 800 34186 856
rect 34354 800 34370 856
rect 34538 800 34554 856
rect 34722 800 34738 856
rect 34906 800 34922 856
rect 35090 800 35106 856
rect 35274 800 35290 856
rect 35458 800 35474 856
rect 35642 800 35658 856
rect 35826 800 35842 856
rect 36010 800 36026 856
rect 36194 800 36210 856
rect 36378 800 36394 856
rect 36562 800 36578 856
rect 36746 800 36762 856
rect 36930 800 36946 856
rect 37114 800 37130 856
rect 37298 800 37314 856
rect 37482 800 37498 856
rect 37666 800 37682 856
rect 37850 800 37866 856
rect 38034 800 38050 856
rect 38218 800 38234 856
rect 38402 800 38418 856
rect 38586 800 38602 856
rect 38770 800 38786 856
rect 38954 800 38970 856
rect 39138 800 39154 856
rect 39322 800 39338 856
rect 39506 800 39522 856
rect 39690 800 39706 856
rect 39874 800 39890 856
rect 40058 800 40074 856
rect 40242 800 40258 856
rect 40426 800 40442 856
rect 40610 800 40626 856
rect 40794 800 40810 856
rect 40978 800 40994 856
rect 41162 800 41178 856
rect 41346 800 41362 856
rect 41530 800 41546 856
rect 41714 800 41730 856
rect 41898 800 41914 856
rect 42082 800 42098 856
rect 42266 800 42282 856
rect 42450 800 42466 856
rect 42634 800 42650 856
rect 42818 800 42834 856
rect 43002 800 43018 856
rect 43186 800 43202 856
rect 43370 800 43386 856
rect 43554 800 43570 856
rect 43738 800 43754 856
rect 43922 800 43938 856
rect 44106 800 44122 856
rect 44290 800 44306 856
rect 44474 800 44490 856
rect 44658 800 44674 856
rect 44842 800 44858 856
rect 45026 800 45042 856
rect 45210 800 45226 856
rect 45394 800 45410 856
rect 45578 800 45594 856
rect 45762 800 45778 856
rect 45946 800 45962 856
rect 46130 800 46146 856
rect 46314 800 46330 856
rect 46498 800 46514 856
rect 46682 800 46698 856
rect 46866 800 46882 856
rect 47050 800 47066 856
rect 47234 800 47250 856
rect 47418 800 47434 856
rect 47602 800 47618 856
rect 47786 800 47802 856
rect 47970 800 47986 856
rect 48154 800 48170 856
rect 48338 800 48354 856
rect 48522 800 48538 856
rect 48706 800 48722 856
rect 48890 800 48906 856
rect 49074 800 49090 856
rect 49258 800 49274 856
rect 49442 800 49458 856
rect 49626 800 49642 856
rect 49810 800 49826 856
rect 49994 800 50010 856
rect 50178 800 50194 856
rect 50362 800 50378 856
rect 50546 800 50562 856
rect 50730 800 50746 856
rect 50914 800 50930 856
rect 51098 800 51114 856
rect 51282 800 51298 856
rect 51466 800 51482 856
rect 51650 800 51666 856
rect 51834 800 51850 856
rect 52018 800 52034 856
rect 52202 800 52218 856
rect 52386 800 52402 856
rect 52570 800 52586 856
rect 52754 800 52770 856
rect 52938 800 52954 856
rect 53122 800 53138 856
rect 53306 800 53322 856
rect 53490 800 53506 856
rect 53674 800 53690 856
rect 53858 800 53874 856
rect 54042 800 54058 856
rect 54226 800 54242 856
rect 54410 800 54426 856
rect 54594 800 54610 856
rect 54778 800 54794 856
rect 54962 800 54978 856
rect 55146 800 55162 856
rect 55330 800 55346 856
rect 55514 800 55530 856
rect 55698 800 55714 856
rect 55882 800 55898 856
rect 56066 800 56082 856
rect 56250 800 56266 856
rect 56434 800 56450 856
rect 56618 800 56634 856
rect 56802 800 56818 856
rect 56986 800 57002 856
rect 57170 800 57186 856
rect 57354 800 57370 856
rect 57538 800 57554 856
rect 57722 800 57738 856
rect 57906 800 57922 856
rect 58090 800 58106 856
rect 58274 800 58290 856
rect 58458 800 58474 856
rect 58642 800 58658 856
rect 58826 800 58842 856
rect 59010 800 59026 856
rect 59194 800 59210 856
rect 59378 800 59394 856
rect 59562 800 59578 856
rect 59746 800 59762 856
rect 59930 800 59946 856
rect 60114 800 60130 856
rect 60298 800 60314 856
rect 60482 800 60498 856
rect 60666 800 60682 856
rect 60850 800 60866 856
rect 61034 800 61050 856
rect 61218 800 61234 856
rect 61402 800 61418 856
rect 61586 800 61602 856
rect 61770 800 61786 856
rect 61954 800 61970 856
rect 62138 800 62154 856
rect 62322 800 62338 856
rect 62506 800 62522 856
rect 62690 800 62706 856
rect 62874 800 62890 856
rect 63058 800 63074 856
rect 63242 800 63258 856
rect 63426 800 63442 856
rect 63610 800 63626 856
rect 63794 800 63810 856
rect 63978 800 63994 856
rect 64162 800 64178 856
rect 64346 800 64362 856
rect 64530 800 64546 856
rect 64714 800 64730 856
rect 64898 800 64914 856
rect 65082 800 65098 856
rect 65266 800 65282 856
rect 65450 800 65466 856
rect 65634 800 65650 856
rect 65818 800 65834 856
rect 66002 800 66018 856
rect 66186 800 66202 856
rect 66370 800 66386 856
rect 66554 800 66570 856
rect 66738 800 66754 856
rect 66922 800 66938 856
rect 67106 800 67122 856
rect 67290 800 67306 856
rect 67474 800 67490 856
rect 67658 800 67674 856
rect 67842 800 67858 856
rect 68026 800 68042 856
rect 68210 800 68226 856
rect 68394 800 68410 856
rect 68578 800 68594 856
rect 68762 800 68778 856
rect 68946 800 68962 856
rect 69130 800 69146 856
rect 69314 800 69330 856
rect 69498 800 69514 856
rect 69682 800 69698 856
rect 69866 800 69882 856
rect 70050 800 70066 856
rect 70234 800 70250 856
rect 70418 800 70434 856
rect 70602 800 70618 856
rect 70786 800 70802 856
rect 70970 800 70986 856
rect 71154 800 71170 856
rect 71338 800 71354 856
rect 71522 800 71538 856
rect 71706 800 71722 856
rect 71890 800 71906 856
rect 72074 800 72090 856
rect 72258 800 72274 856
rect 72442 800 72458 856
rect 72626 800 72642 856
rect 72810 800 72826 856
rect 72994 800 73010 856
rect 73178 800 73194 856
rect 73362 800 73378 856
rect 73546 800 73562 856
rect 73730 800 73746 856
rect 73914 800 73930 856
rect 74098 800 74114 856
rect 74282 800 74298 856
rect 74466 800 74482 856
rect 74650 800 74666 856
rect 74834 800 74850 856
rect 75018 800 75034 856
rect 75202 800 75218 856
rect 75386 800 75402 856
rect 75570 800 75586 856
rect 75754 800 75770 856
rect 75938 800 75954 856
rect 76122 800 76138 856
rect 76306 800 76322 856
rect 76490 800 76506 856
rect 76674 800 76690 856
rect 76858 800 76874 856
rect 77042 800 77058 856
rect 77226 800 77242 856
rect 77410 800 77426 856
rect 77594 800 77610 856
rect 77778 800 77794 856
rect 77962 800 77978 856
rect 78146 800 78162 856
rect 78330 800 78346 856
rect 78514 800 78530 856
rect 78698 800 78714 856
rect 78882 800 78898 856
rect 79066 800 79082 856
rect 79250 800 79266 856
rect 79434 800 79450 856
rect 79618 800 79634 856
rect 79802 800 79818 856
rect 79986 800 80002 856
rect 80170 800 80186 856
rect 80354 800 80370 856
rect 80538 800 80554 856
rect 80722 800 80738 856
rect 80906 800 80922 856
rect 81090 800 81106 856
rect 81274 800 81290 856
rect 81458 800 81474 856
rect 81642 800 81658 856
rect 81826 800 81842 856
rect 82010 800 82026 856
rect 82194 800 82210 856
rect 82378 800 82394 856
rect 82562 800 82578 856
rect 82746 800 82762 856
rect 82930 800 82946 856
rect 83114 800 83130 856
rect 83298 800 83314 856
rect 83482 800 83498 856
rect 83666 800 83682 856
rect 83850 800 83866 856
rect 84034 800 84050 856
rect 84218 800 84234 856
rect 84402 800 84418 856
rect 84586 800 84602 856
rect 84770 800 84786 856
rect 84954 800 84970 856
rect 85138 800 85154 856
rect 85322 800 85338 856
rect 85506 800 85522 856
rect 85690 800 85706 856
rect 85874 800 85890 856
rect 86058 800 86074 856
rect 86242 800 86258 856
rect 86426 800 86442 856
rect 86610 800 86626 856
rect 86794 800 86810 856
rect 86978 800 86994 856
rect 87162 800 87178 856
rect 87346 800 87362 856
rect 87530 800 87546 856
rect 87714 800 87730 856
rect 87898 800 87914 856
rect 88082 800 88098 856
rect 88266 800 88282 856
rect 88450 800 88466 856
rect 88634 800 88650 856
rect 88818 800 88834 856
rect 89002 800 89018 856
rect 89186 800 89202 856
rect 89370 800 89386 856
rect 89554 800 89570 856
rect 89738 800 89754 856
rect 89922 800 89938 856
rect 90106 800 90122 856
rect 90290 800 90306 856
rect 90474 800 90490 856
rect 90658 800 90674 856
rect 90842 800 90858 856
rect 91026 800 91042 856
rect 91210 800 91226 856
rect 91394 800 91410 856
rect 91578 800 91594 856
rect 91762 800 91778 856
rect 91946 800 91962 856
rect 92130 800 92146 856
rect 92314 800 92330 856
rect 92498 800 92514 856
rect 92682 800 92698 856
rect 92866 800 92882 856
rect 93050 800 93066 856
rect 93234 800 93250 856
rect 93418 800 93434 856
rect 93602 800 93618 856
rect 93786 800 93802 856
rect 93970 800 93986 856
rect 94154 800 94170 856
rect 94338 800 94354 856
rect 94522 800 94538 856
rect 94706 800 94722 856
rect 94890 800 94906 856
rect 95074 800 95090 856
rect 95258 800 95274 856
rect 95442 800 95458 856
rect 95626 800 95642 856
rect 95810 800 95826 856
rect 95994 800 96010 856
rect 96178 800 96194 856
rect 96362 800 96378 856
rect 96546 800 96562 856
rect 96730 800 96746 856
rect 96914 800 96930 856
rect 97098 800 97114 856
rect 97282 800 97298 856
rect 97466 800 97482 856
rect 97650 800 97666 856
rect 97834 800 97850 856
rect 98018 800 98034 856
rect 98202 800 98218 856
rect 98386 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98770 856
rect 98938 800 98954 856
rect 99122 800 99138 856
rect 99306 800 99322 856
rect 99490 800 99506 856
rect 99674 800 99690 856
rect 99858 800 99874 856
rect 100042 800 100058 856
rect 100226 800 100242 856
rect 100410 800 100426 856
rect 100594 800 100610 856
rect 100778 800 100794 856
rect 100962 800 100978 856
rect 101146 800 101162 856
rect 101330 800 101346 856
rect 101514 800 101530 856
rect 101698 800 101714 856
rect 101882 800 101898 856
rect 102066 800 102082 856
rect 102250 800 102266 856
rect 102434 800 102450 856
rect 102618 800 102634 856
rect 102802 800 102818 856
rect 102986 800 103002 856
rect 103170 800 103186 856
rect 103354 800 103370 856
rect 103538 800 103554 856
rect 103722 800 103738 856
rect 103906 800 103922 856
rect 104090 800 104106 856
rect 104274 800 104290 856
rect 104458 800 104474 856
rect 104642 800 104658 856
rect 104826 800 104842 856
rect 105010 800 105026 856
rect 105194 800 105210 856
rect 105378 800 105394 856
rect 105562 800 105578 856
rect 105746 800 105762 856
rect 105930 800 105946 856
rect 106114 800 106130 856
rect 106298 800 106314 856
rect 106482 800 106498 856
rect 106666 800 106682 856
rect 106850 800 106866 856
rect 107034 800 107050 856
rect 107218 800 107234 856
rect 107402 800 107418 856
rect 107586 800 107602 856
rect 107770 800 107786 856
rect 107954 800 107970 856
rect 108138 800 108154 856
rect 108322 800 108338 856
rect 108506 800 108522 856
rect 108690 800 108706 856
rect 108874 800 108890 856
rect 109058 800 109074 856
rect 109242 800 109258 856
rect 109426 800 109442 856
rect 109610 800 109626 856
rect 109794 800 109810 856
rect 109978 800 109994 856
rect 110162 800 110178 856
rect 110346 800 129240 856
<< metal3 >>
rect 129284 128936 130084 129056
rect 0 126760 800 126880
rect 0 124584 800 124704
rect 129284 124584 130084 124704
rect 0 122408 800 122528
rect 0 120232 800 120352
rect 129284 120232 130084 120352
rect 0 118056 800 118176
rect 0 115880 800 116000
rect 129284 115880 130084 116000
rect 0 113704 800 113824
rect 0 111528 800 111648
rect 129284 111528 130084 111648
rect 0 109352 800 109472
rect 0 107176 800 107296
rect 129284 107176 130084 107296
rect 0 105000 800 105120
rect 0 102824 800 102944
rect 129284 102824 130084 102944
rect 0 100648 800 100768
rect 0 98472 800 98592
rect 129284 98472 130084 98592
rect 0 96296 800 96416
rect 0 94120 800 94240
rect 129284 94120 130084 94240
rect 0 91944 800 92064
rect 0 89768 800 89888
rect 129284 89768 130084 89888
rect 0 87592 800 87712
rect 0 85416 800 85536
rect 129284 85416 130084 85536
rect 0 83240 800 83360
rect 0 81064 800 81184
rect 129284 81064 130084 81184
rect 0 78888 800 79008
rect 0 76712 800 76832
rect 129284 76712 130084 76832
rect 0 74536 800 74656
rect 0 72360 800 72480
rect 129284 72360 130084 72480
rect 0 70184 800 70304
rect 0 68008 800 68128
rect 129284 68008 130084 68128
rect 0 65832 800 65952
rect 0 63656 800 63776
rect 129284 63656 130084 63776
rect 0 61480 800 61600
rect 0 59304 800 59424
rect 129284 59304 130084 59424
rect 0 57128 800 57248
rect 0 54952 800 55072
rect 129284 54952 130084 55072
rect 0 52776 800 52896
rect 0 50600 800 50720
rect 129284 50600 130084 50720
rect 0 48424 800 48544
rect 0 46248 800 46368
rect 129284 46248 130084 46368
rect 0 44072 800 44192
rect 0 41896 800 42016
rect 129284 41896 130084 42016
rect 0 39720 800 39840
rect 0 37544 800 37664
rect 129284 37544 130084 37664
rect 0 35368 800 35488
rect 0 33192 800 33312
rect 129284 33192 130084 33312
rect 0 31016 800 31136
rect 0 28840 800 28960
rect 129284 28840 130084 28960
rect 0 26664 800 26784
rect 0 24488 800 24608
rect 129284 24488 130084 24608
rect 0 22312 800 22432
rect 0 20136 800 20256
rect 129284 20136 130084 20256
rect 0 17960 800 18080
rect 0 15784 800 15904
rect 129284 15784 130084 15904
rect 0 13608 800 13728
rect 0 11432 800 11552
rect 129284 11432 130084 11552
rect 0 9256 800 9376
rect 0 7080 800 7200
rect 129284 7080 130084 7200
rect 0 4904 800 5024
rect 129284 2728 130084 2848
<< obsm3 >>
rect 798 129136 129284 130049
rect 798 128856 129204 129136
rect 798 126960 129284 128856
rect 880 126680 129284 126960
rect 798 124784 129284 126680
rect 880 124504 129204 124784
rect 798 122608 129284 124504
rect 880 122328 129284 122608
rect 798 120432 129284 122328
rect 880 120152 129204 120432
rect 798 118256 129284 120152
rect 880 117976 129284 118256
rect 798 116080 129284 117976
rect 880 115800 129204 116080
rect 798 113904 129284 115800
rect 880 113624 129284 113904
rect 798 111728 129284 113624
rect 880 111448 129204 111728
rect 798 109552 129284 111448
rect 880 109272 129284 109552
rect 798 107376 129284 109272
rect 880 107096 129204 107376
rect 798 105200 129284 107096
rect 880 104920 129284 105200
rect 798 103024 129284 104920
rect 880 102744 129204 103024
rect 798 100848 129284 102744
rect 880 100568 129284 100848
rect 798 98672 129284 100568
rect 880 98392 129204 98672
rect 798 96496 129284 98392
rect 880 96216 129284 96496
rect 798 94320 129284 96216
rect 880 94040 129204 94320
rect 798 92144 129284 94040
rect 880 91864 129284 92144
rect 798 89968 129284 91864
rect 880 89688 129204 89968
rect 798 87792 129284 89688
rect 880 87512 129284 87792
rect 798 85616 129284 87512
rect 880 85336 129204 85616
rect 798 83440 129284 85336
rect 880 83160 129284 83440
rect 798 81264 129284 83160
rect 880 80984 129204 81264
rect 798 79088 129284 80984
rect 880 78808 129284 79088
rect 798 76912 129284 78808
rect 880 76632 129204 76912
rect 798 74736 129284 76632
rect 880 74456 129284 74736
rect 798 72560 129284 74456
rect 880 72280 129204 72560
rect 798 70384 129284 72280
rect 880 70104 129284 70384
rect 798 68208 129284 70104
rect 880 67928 129204 68208
rect 798 66032 129284 67928
rect 880 65752 129284 66032
rect 798 63856 129284 65752
rect 880 63576 129204 63856
rect 798 61680 129284 63576
rect 880 61400 129284 61680
rect 798 59504 129284 61400
rect 880 59224 129204 59504
rect 798 57328 129284 59224
rect 880 57048 129284 57328
rect 798 55152 129284 57048
rect 880 54872 129204 55152
rect 798 52976 129284 54872
rect 880 52696 129284 52976
rect 798 50800 129284 52696
rect 880 50520 129204 50800
rect 798 48624 129284 50520
rect 880 48344 129284 48624
rect 798 46448 129284 48344
rect 880 46168 129204 46448
rect 798 44272 129284 46168
rect 880 43992 129284 44272
rect 798 42096 129284 43992
rect 880 41816 129204 42096
rect 798 39920 129284 41816
rect 880 39640 129284 39920
rect 798 37744 129284 39640
rect 880 37464 129204 37744
rect 798 35568 129284 37464
rect 880 35288 129284 35568
rect 798 33392 129284 35288
rect 880 33112 129204 33392
rect 798 31216 129284 33112
rect 880 30936 129284 31216
rect 798 29040 129284 30936
rect 880 28760 129204 29040
rect 798 26864 129284 28760
rect 880 26584 129284 26864
rect 798 24688 129284 26584
rect 880 24408 129204 24688
rect 798 22512 129284 24408
rect 880 22232 129284 22512
rect 798 20336 129284 22232
rect 880 20056 129204 20336
rect 798 18160 129284 20056
rect 880 17880 129284 18160
rect 798 15984 129284 17880
rect 880 15704 129204 15984
rect 798 13808 129284 15704
rect 880 13528 129284 13808
rect 798 11632 129284 13528
rect 880 11352 129204 11632
rect 798 9456 129284 11352
rect 880 9176 129284 9456
rect 798 7280 129284 9176
rect 880 7000 129204 7280
rect 798 5104 129284 7000
rect 880 4824 129284 5104
rect 798 2928 129284 4824
rect 798 2648 129204 2928
rect 798 1803 129284 2648
<< metal4 >>
rect 3748 2128 4988 130064
rect 13748 2128 14988 130064
rect 23748 2128 24988 130064
rect 33748 2128 34988 130064
rect 43748 2128 44988 130064
rect 53748 2128 54988 130064
rect 63748 2128 64988 130064
rect 73748 2128 74988 130064
rect 83748 2128 84988 130064
rect 93748 2128 94988 130064
rect 103748 2128 104988 130064
rect 113748 2128 114988 130064
rect 123748 2128 124988 130064
<< obsm4 >>
rect 11099 2048 13668 129709
rect 15068 2048 23668 129709
rect 25068 2048 33668 129709
rect 35068 2048 43668 129709
rect 45068 2048 53668 129709
rect 55068 2048 63668 129709
rect 65068 2048 73668 129709
rect 75068 2048 83668 129709
rect 85068 2048 93668 129709
rect 95068 2048 103668 129709
rect 105068 2048 113668 129709
rect 115068 2048 123668 129709
rect 125068 2048 128189 129709
rect 11099 1803 128189 2048
<< labels >>
rlabel metal3 s 129284 2728 130084 2848 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 127162 131428 127218 132228 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 112810 131428 112866 132228 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 98458 131428 98514 132228 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 84106 131428 84162 132228 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 69754 131428 69810 132228 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 55402 131428 55458 132228 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 41050 131428 41106 132228 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 26698 131428 26754 132228 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 12346 131428 12402 132228 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 126760 800 126880 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 129284 15784 130084 15904 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 120232 800 120352 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 113704 800 113824 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 129284 28840 130084 28960 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 129284 41896 130084 42016 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 129284 54952 130084 55072 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 129284 68008 130084 68128 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 129284 81064 130084 81184 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 129284 94120 130084 94240 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 129284 107176 130084 107296 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 129284 120232 130084 120352 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 129284 11432 130084 11552 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 117594 131428 117650 132228 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 103242 131428 103298 132228 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 88890 131428 88946 132228 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 74538 131428 74594 132228 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 60186 131428 60242 132228 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 45834 131428 45890 132228 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 31482 131428 31538 132228 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 17130 131428 17186 132228 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 2778 131428 2834 132228 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 129284 24488 130084 24608 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 102824 800 102944 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 0 96296 800 96416 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 76712 800 76832 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 70184 800 70304 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 129284 37544 130084 37664 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 50600 800 50720 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 129284 50600 130084 50720 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 129284 63656 130084 63776 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 129284 76712 130084 76832 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 129284 89768 130084 89888 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 129284 102824 130084 102944 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 129284 115880 130084 116000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 129284 128936 130084 129056 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 129284 7080 130084 7200 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 122378 131428 122434 132228 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 108026 131428 108082 132228 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 93674 131428 93730 132228 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 79322 131428 79378 132228 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 64970 131428 65026 132228 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 50618 131428 50674 132228 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 36266 131428 36322 132228 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 21914 131428 21970 132228 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 7562 131428 7618 132228 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 129284 20136 130084 20256 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 0 105000 800 105120 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 0 98472 800 98592 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 91944 800 92064 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 72360 800 72480 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 65832 800 65952 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 129284 33192 130084 33312 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 129284 46248 130084 46368 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 129284 59304 130084 59424 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 129284 72360 130084 72480 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 129284 85416 130084 85536 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 129284 98472 130084 98592 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 129284 111528 130084 111648 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 129284 124584 130084 124704 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 99562 0 99618 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 108946 0 109002 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 87970 0 88026 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 3748 2128 4988 130064 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 23748 2128 24988 130064 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 43748 2128 44988 130064 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 63748 2128 64988 130064 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 83748 2128 84988 130064 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 103748 2128 104988 130064 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 123748 2128 124988 130064 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 13748 2128 14988 130064 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 33748 2128 34988 130064 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 53748 2128 54988 130064 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 73748 2128 74988 130064 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 93748 2128 94988 130064 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 113748 2128 114988 130064 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 19706 0 19762 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 130084 132228
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 67997102
string GDS_FILE /home/ejjimenezu/Repos/caravel_simple_fpu/openlane/fpu/runs/24_12_05_06_12/results/signoff/fpu.magic.gds
string GDS_START 1073570
<< end >>

